/**
 * Copyright (C) 2020  AGH University of Science and Technology
 *
 * This program is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with this program.  If not, see <https://www.gnu.org/licenses/>.
 */

module spi_mem (
    output logic [31:0] rdata,
    input logic [31:0] addr
);

/**
 * Module internal logic
 */

always_comb begin
    case (addr[13:2])
           0:    rdata = 32'h08c0006f;
           1:    rdata = 32'h0880006f;
           2:    rdata = 32'h0840006f;
           3:    rdata = 32'h0800006f;
           4:    rdata = 32'h07c0006f;
           5:    rdata = 32'h0780006f;
           6:    rdata = 32'h0740006f;
           7:    rdata = 32'h0700006f;
           8:    rdata = 32'h06c0006f;
           9:    rdata = 32'h0680006f;
          10:    rdata = 32'h0640006f;
          11:    rdata = 32'h0600006f;
          12:    rdata = 32'h05c0006f;
          13:    rdata = 32'h0580006f;
          14:    rdata = 32'h0540006f;
          15:    rdata = 32'h0500006f;
          16:    rdata = 32'h1e40106f;
          17:    rdata = 32'h2320106f;
          18:    rdata = 32'h0440006f;
          19:    rdata = 32'h0400006f;
          20:    rdata = 32'h03c0006f;
          21:    rdata = 32'h0380006f;
          22:    rdata = 32'h0340006f;
          23:    rdata = 32'h0300006f;
          24:    rdata = 32'h02c0006f;
          25:    rdata = 32'h0280006f;
          26:    rdata = 32'h0240006f;
          27:    rdata = 32'h0200006f;
          28:    rdata = 32'h01c0006f;
          29:    rdata = 32'h0180006f;
          30:    rdata = 32'h0140006f;
          31:    rdata = 32'h0100006f;
          32:    rdata = 32'h0100006f;
          33:    rdata = 32'h0080006f;
          34:    rdata = 32'h0040006f;
          35:    rdata = 32'h0000006f;
          36:    rdata = 32'h00000093;
          37:    rdata = 32'h00000113;
          38:    rdata = 32'h00000193;
          39:    rdata = 32'h00000213;
          40:    rdata = 32'h00000293;
          41:    rdata = 32'h00000313;
          42:    rdata = 32'h00000393;
          43:    rdata = 32'h00000413;
          44:    rdata = 32'h00000493;
          45:    rdata = 32'h00000513;
          46:    rdata = 32'h00000593;
          47:    rdata = 32'h00000613;
          48:    rdata = 32'h00000693;
          49:    rdata = 32'h00000713;
          50:    rdata = 32'h00000793;
          51:    rdata = 32'h00000813;
          52:    rdata = 32'h00000893;
          53:    rdata = 32'h00000913;
          54:    rdata = 32'h00000993;
          55:    rdata = 32'h00000a13;
          56:    rdata = 32'h00000a93;
          57:    rdata = 32'h00000b13;
          58:    rdata = 32'h00000b93;
          59:    rdata = 32'h00000c13;
          60:    rdata = 32'h00000c93;
          61:    rdata = 32'h00000d13;
          62:    rdata = 32'h00000d93;
          63:    rdata = 32'h00000e13;
          64:    rdata = 32'h00000e93;
          65:    rdata = 32'h00000f13;
          66:    rdata = 32'h00000f93;
          67:    rdata = 32'h000f4117;
          68:    rdata = 32'hef410113;
          69:    rdata = 32'h000f0297;
          70:    rdata = 32'heec28293;
          71:    rdata = 32'h000f0317;
          72:    rdata = 32'hf7030313;
          73:    rdata = 32'h0062d863;
          74:    rdata = 32'h0002a023;
          75:    rdata = 32'h00428293;
          76:    rdata = 32'hfe535ce3;
          77:    rdata = 32'h00002297;
          78:    rdata = 32'hce428293;
          79:    rdata = 32'h000f0317;
          80:    rdata = 32'hec430313;
          81:    rdata = 32'h000f0397;
          82:    rdata = 32'hebc38393;
          83:    rdata = 32'h00735c63;
          84:    rdata = 32'h0002ae03;
          85:    rdata = 32'h01c32023;
          86:    rdata = 32'h00428293;
          87:    rdata = 32'h00430313;
          88:    rdata = 32'hfe7348e3;
          89:    rdata = 32'h00001297;
          90:    rdata = 32'h78428293;
          91:    rdata = 32'h00001317;
          92:    rdata = 32'h79030313;
          93:    rdata = 32'h0062da63;
          94:    rdata = 32'h0002a783;
          95:    rdata = 32'h000780e7;
          96:    rdata = 32'h00428293;
          97:    rdata = 32'hfe62cae3;
          98:    rdata = 32'h00000513;
          99:    rdata = 32'h00000593;
         100:    rdata = 32'h6c0010ef;
         101:    rdata = 32'h25971141;
         102:    rdata = 32'h85930000;
         103:    rdata = 32'h05178125;
         104:    rdata = 32'h0513000f;
         105:    rdata = 32'hc606eda5;
         106:    rdata = 32'h787000ef;
         107:    rdata = 32'h051740b2;
         108:    rdata = 32'h0513000f;
         109:    rdata = 32'h0141ea25;
         110:    rdata = 32'h3a80106f;
         111:    rdata = 32'h00001597;
         112:    rdata = 32'h7f858593;
         113:    rdata = 32'h000f0517;
         114:    rdata = 32'heb450513;
         115:    rdata = 32'h7630006f;
         116:    rdata = 32'h00002597;
         117:    rdata = 32'ha0058593;
         118:    rdata = 32'h000f0517;
         119:    rdata = 32'hea050513;
         120:    rdata = 32'h74f0006f;
         121:    rdata = 32'h00002597;
         122:    rdata = 32'ha0c58593;
         123:    rdata = 32'h000f0517;
         124:    rdata = 32'he8c50513;
         125:    rdata = 32'h73b0006f;
         126:    rdata = 32'h114141d8;
         127:    rdata = 32'hc422c606;
         128:    rdata = 32'hc04ac226;
         129:    rdata = 32'hc4634785;
         130:    rdata = 32'h259702e7;
         131:    rdata = 32'h85930000;
         132:    rdata = 32'h05179ee5;
         133:    rdata = 32'h0513000f;
         134:    rdata = 32'h00efe665;
         135:    rdata = 32'h44057150;
         136:    rdata = 32'h852240b2;
         137:    rdata = 32'h44924422;
         138:    rdata = 32'h01414902;
         139:    rdata = 32'h45808082;
         140:    rdata = 32'h146384ae;
         141:    rdata = 32'h519c00f4;
         142:    rdata = 32'h2597c791;
         143:    rdata = 32'h85930000;
         144:    rdata = 32'hbfc19da5;
         145:    rdata = 32'h02458913;
         146:    rdata = 32'h2597854a;
         147:    rdata = 32'h85930000;
         148:    rdata = 32'h00ef9ee5;
         149:    rdata = 32'hc50d4750;
         150:    rdata = 32'h00002597;
         151:    rdata = 32'h9e458593;
         152:    rdata = 32'h00ef854a;
         153:    rdata = 32'hcd014650;
         154:    rdata = 32'h00002597;
         155:    rdata = 32'h9d858593;
         156:    rdata = 32'h000f0517;
         157:    rdata = 32'he0850513;
         158:    rdata = 32'h6b7000ef;
         159:    rdata = 32'h4401b755;
         160:    rdata = 32'h00c4c583;
         161:    rdata = 32'h05178622;
         162:    rdata = 32'h0513000f;
         163:    rdata = 32'h10efd7a5;
         164:    rdata = 32'h440106e0;
         165:    rdata = 32'h41dcb771;
         166:    rdata = 32'hc6061141;
         167:    rdata = 32'h02f04063;
         168:    rdata = 32'h00002597;
         169:    rdata = 32'h9bc58593;
         170:    rdata = 32'h000f0517;
         171:    rdata = 32'hdd050513;
         172:    rdata = 32'h67f000ef;
         173:    rdata = 32'h40b24505;
         174:    rdata = 32'h80820141;
         175:    rdata = 32'h47854598;
         176:    rdata = 32'h00f70763;
         177:    rdata = 32'h00002597;
         178:    rdata = 32'h9b458593;
         179:    rdata = 32'hc583bff1;
         180:    rdata = 32'h051700c5;
         181:    rdata = 32'h0513000f;
         182:    rdata = 32'h10efd2e5;
         183:    rdata = 32'h25970380;
         184:    rdata = 32'h85930000;
         185:    rdata = 32'hc50995e5;
         186:    rdata = 32'h00002597;
         187:    rdata = 32'h95058593;
         188:    rdata = 32'h000f0517;
         189:    rdata = 32'hd8850513;
         190:    rdata = 32'h637000ef;
         191:    rdata = 32'h00002597;
         192:    rdata = 32'h99858593;
         193:    rdata = 32'h62b000ef;
         194:    rdata = 32'hb7754501;
         195:    rdata = 32'h114141dc;
         196:    rdata = 32'h4705c606;
         197:    rdata = 32'h02f74063;
         198:    rdata = 32'h00002597;
         199:    rdata = 32'h8e058593;
         200:    rdata = 32'h000f0517;
         201:    rdata = 32'hd5850513;
         202:    rdata = 32'h607000ef;
         203:    rdata = 32'h40b24505;
         204:    rdata = 32'h80820141;
         205:    rdata = 32'h9563459c;
         206:    rdata = 32'h519800e7;
         207:    rdata = 32'h00f70763;
         208:    rdata = 32'h00002597;
         209:    rdata = 32'h8d458593;
         210:    rdata = 32'h51d0bfe1;
         211:    rdata = 32'h00c5c583;
         212:    rdata = 32'h000f0517;
         213:    rdata = 32'hcb050513;
         214:    rdata = 32'h00c03633;
         215:    rdata = 32'h7eb000ef;
         216:    rdata = 32'hb7f14501;
         217:    rdata = 32'h110141dc;
         218:    rdata = 32'h4063ce06;
         219:    rdata = 32'h259702f0;
         220:    rdata = 32'h85930000;
         221:    rdata = 32'h05178ee5;
         222:    rdata = 32'h0513000f;
         223:    rdata = 32'h00efd025;
         224:    rdata = 32'h45055b10;
         225:    rdata = 32'h610540f2;
         226:    rdata = 32'h45988082;
         227:    rdata = 32'h07634785;
         228:    rdata = 32'h259700f7;
         229:    rdata = 32'h85930000;
         230:    rdata = 32'hbff18e65;
         231:    rdata = 32'h00c5c583;
         232:    rdata = 32'h000f0517;
         233:    rdata = 32'hc6050513;
         234:    rdata = 32'h77d000ef;
         235:    rdata = 32'h006cc62a;
         236:    rdata = 32'h000f0517;
         237:    rdata = 32'hcc850513;
         238:    rdata = 32'h593000ef;
         239:    rdata = 32'h00002597;
         240:    rdata = 32'h8d858593;
         241:    rdata = 32'h56b000ef;
         242:    rdata = 32'hbf6d4501;
         243:    rdata = 32'h114141dc;
         244:    rdata = 32'hc422c606;
         245:    rdata = 32'h02f04163;
         246:    rdata = 32'h00002597;
         247:    rdata = 32'h88458593;
         248:    rdata = 32'h000f0517;
         249:    rdata = 32'hc9850513;
         250:    rdata = 32'h547000ef;
         251:    rdata = 32'h40b24505;
         252:    rdata = 32'h01414422;
         253:    rdata = 32'h45988082;
         254:    rdata = 32'h842e4785;
         255:    rdata = 32'h00f70763;
         256:    rdata = 32'h00002597;
         257:    rdata = 32'h87858593;
         258:    rdata = 32'h45dcbfe1;
         259:    rdata = 32'h04f05363;
         260:    rdata = 32'h00000597;
         261:    rdata = 32'hd8458593;
         262:    rdata = 32'h000f0517;
         263:    rdata = 32'hc6450513;
         264:    rdata = 32'h5eb000ef;
         265:    rdata = 32'h6731445c;
         266:    rdata = 32'h35070713;
         267:    rdata = 32'h02e787b3;
         268:    rdata = 32'h000f0517;
         269:    rdata = 32'hc2050513;
         270:    rdata = 32'h17fd4558;
         271:    rdata = 32'h10efc31c;
         272:    rdata = 32'h051710c0;
         273:    rdata = 32'h0513000f;
         274:    rdata = 32'h00efc3a5;
         275:    rdata = 32'h450159f0;
         276:    rdata = 32'h0517bf79;
         277:    rdata = 32'h0513000f;
         278:    rdata = 32'h10efbfe5;
         279:    rdata = 32'h05170fc0;
         280:    rdata = 32'h0513000f;
         281:    rdata = 32'h00efc1e5;
         282:    rdata = 32'hb7d55b10;
         283:    rdata = 32'hce061101;
         284:    rdata = 32'hca26cc22;
         285:    rdata = 32'h81010113;
         286:    rdata = 32'h04000613;
         287:    rdata = 32'h850a4581;
         288:    rdata = 32'h2f4010ef;
         289:    rdata = 32'h0517858a;
         290:    rdata = 32'h0513000f;
         291:    rdata = 32'h00efb9e5;
         292:    rdata = 32'h051774d0;
         293:    rdata = 32'h0513000f;
         294:    rdata = 32'h00efbea5;
         295:    rdata = 32'h842a5330;
         296:    rdata = 32'h000f0597;
         297:    rdata = 32'hbd458593;
         298:    rdata = 32'h2b4d850a;
         299:    rdata = 32'h000f0517;
         300:    rdata = 32'hbd050513;
         301:    rdata = 32'h519000ef;
         302:    rdata = 32'h408505b3;
         303:    rdata = 32'h00001517;
         304:    rdata = 32'h7dc50513;
         305:    rdata = 32'h840a2935;
         306:    rdata = 32'h55030084;
         307:    rdata = 32'h04097c04;
         308:    rdata = 32'h1ce32ee1;
         309:    rdata = 32'h0113fe94;
         310:    rdata = 32'h40f27f01;
         311:    rdata = 32'h44d24462;
         312:    rdata = 32'h80826105;
         313:    rdata = 32'h0593715d;
         314:    rdata = 32'h05170400;
         315:    rdata = 32'h0513000f;
         316:    rdata = 32'hc686b3a5;
         317:    rdata = 32'h00efc4a2;
         318:    rdata = 32'h06137130;
         319:    rdata = 32'h45810400;
         320:    rdata = 32'h10ef850a;
         321:    rdata = 32'h858a2720;
         322:    rdata = 32'h000f0517;
         323:    rdata = 32'hb1c50513;
         324:    rdata = 32'h6cb000ef;
         325:    rdata = 32'h000f0517;
         326:    rdata = 32'hb6850513;
         327:    rdata = 32'h4b1000ef;
         328:    rdata = 32'h0517842a;
         329:    rdata = 32'h0513000f;
         330:    rdata = 32'h00efb525;
         331:    rdata = 32'h05176980;
         332:    rdata = 32'h0513000f;
         333:    rdata = 32'h00efb4e5;
         334:    rdata = 32'h04334970;
         335:    rdata = 32'h15974085;
         336:    rdata = 32'h85930000;
         337:    rdata = 32'h051776a5;
         338:    rdata = 32'h0513000f;
         339:    rdata = 32'h00efb325;
         340:    rdata = 32'h85a23e10;
         341:    rdata = 32'h40b64426;
         342:    rdata = 32'h00001517;
         343:    rdata = 32'h76c50513;
         344:    rdata = 32'hae796161;
         345:    rdata = 32'h2c23712d;
         346:    rdata = 32'h2a231081;
         347:    rdata = 32'h28231091;
         348:    rdata = 32'h26231121;
         349:    rdata = 32'h24231131;
         350:    rdata = 32'h22231141;
         351:    rdata = 32'h20231151;
         352:    rdata = 32'h2e231161;
         353:    rdata = 32'h842a1011;
         354:    rdata = 32'h00001a97;
         355:    rdata = 32'h750a8a93;
         356:    rdata = 32'h000f0497;
         357:    rdata = 32'hae848493;
         358:    rdata = 32'h19174a29;
         359:    rdata = 32'h09130000;
         360:    rdata = 32'h19973629;
         361:    rdata = 32'h89930000;
         362:    rdata = 32'h1b1778e9;
         363:    rdata = 32'h0b130000;
         364:    rdata = 32'h85d6732b;
         365:    rdata = 32'h00ef8526;
         366:    rdata = 32'h004c3790;
         367:    rdata = 32'h00ef8526;
         368:    rdata = 32'h00503350;
         369:    rdata = 32'h10a885a2;
         370:    rdata = 32'h57a62c99;
         371:    rdata = 32'hfefa63e3;
         372:    rdata = 32'h97ca078a;
         373:    rdata = 32'h97ca439c;
         374:    rdata = 32'h85228782;
         375:    rdata = 32'hbfd136c5;
         376:    rdata = 32'h36fd8522;
         377:    rdata = 32'h8522b7f9;
         378:    rdata = 32'hb7e13ef5;
         379:    rdata = 32'h852210ac;
         380:    rdata = 32'hd1613121;
         381:    rdata = 32'h852685ce;
         382:    rdata = 32'h10aca091;
         383:    rdata = 32'h39618522;
         384:    rdata = 32'h10acbfcd;
         385:    rdata = 32'h33198522;
         386:    rdata = 32'h10acb7ed;
         387:    rdata = 32'h3b998522;
         388:    rdata = 32'h10acb7cd;
         389:    rdata = 32'h3b5d8522;
         390:    rdata = 32'h8522bfe9;
         391:    rdata = 32'hbf513d81;
         392:    rdata = 32'h35c98522;
         393:    rdata = 32'h85dab779;
         394:    rdata = 32'h00ef8526;
         395:    rdata = 32'h004c3050;
         396:    rdata = 32'h2e3000ef;
         397:    rdata = 32'h00001597;
         398:    rdata = 32'h6c858593;
         399:    rdata = 32'h2f3000ef;
         400:    rdata = 32'h852ebf8d;
         401:    rdata = 32'h02000713;
         402:    rdata = 32'h00054783;
         403:    rdata = 32'h9563c789;
         404:    rdata = 32'h050500e7;
         405:    rdata = 32'h4501bfd5;
         406:    rdata = 32'h47838082;
         407:    rdata = 32'hf7130006;
         408:    rdata = 32'hc7110df7;
         409:    rdata = 32'h06050585;
         410:    rdata = 32'hfef58fa3;
         411:    rdata = 32'h8023b7fd;
         412:    rdata = 32'h80820005;
         413:    rdata = 32'h0005c783;
         414:    rdata = 32'h0df7f793;
         415:    rdata = 32'h0585c399;
         416:    rdata = 32'h8513bfd5;
         417:    rdata = 32'h8082fff5;
         418:    rdata = 32'hcc221101;
         419:    rdata = 32'hc452c84a;
         420:    rdata = 32'hc05ac256;
         421:    rdata = 32'hca26ce06;
         422:    rdata = 32'h892ac64e;
         423:    rdata = 32'h4b158432;
         424:    rdata = 32'h00860a13;
         425:    rdata = 32'h40444ae1;
         426:    rdata = 32'h029b4663;
         427:    rdata = 32'h3f51854a;
         428:    rdata = 32'hc10d89aa;
         429:    rdata = 32'h035485b3;
         430:    rdata = 32'h854a862a;
         431:    rdata = 32'h95d20591;
         432:    rdata = 32'h85ce3f69;
         433:    rdata = 32'h377d854a;
         434:    rdata = 32'h0593405c;
         435:    rdata = 32'h07850015;
         436:    rdata = 32'hbfd1c05c;
         437:    rdata = 32'h446240f2;
         438:    rdata = 32'h494244d2;
         439:    rdata = 32'h4a2249b2;
         440:    rdata = 32'h4b024a92;
         441:    rdata = 32'h80826105;
         442:    rdata = 32'hc2261141;
         443:    rdata = 32'h00c58493;
         444:    rdata = 32'h8526c422;
         445:    rdata = 32'h1597842e;
         446:    rdata = 32'h85930000;
         447:    rdata = 32'hc6066525;
         448:    rdata = 32'h7c6000ef;
         449:    rdata = 32'h2023e919;
         450:    rdata = 32'h405c0004;
         451:    rdata = 32'h449240b2;
         452:    rdata = 32'hc05c17fd;
         453:    rdata = 32'h01414422;
         454:    rdata = 32'h15978082;
         455:    rdata = 32'h85930000;
         456:    rdata = 32'h85266365;
         457:    rdata = 32'h7a2000ef;
         458:    rdata = 32'hc9514785;
         459:    rdata = 32'h00001597;
         460:    rdata = 32'h62c58593;
         461:    rdata = 32'h00ef8526;
         462:    rdata = 32'h47897900;
         463:    rdata = 32'h1597c149;
         464:    rdata = 32'h85930000;
         465:    rdata = 32'h85266225;
         466:    rdata = 32'h77e000ef;
         467:    rdata = 32'hc925478d;
         468:    rdata = 32'h00001597;
         469:    rdata = 32'h62458593;
         470:    rdata = 32'h00ef8526;
         471:    rdata = 32'h479176c0;
         472:    rdata = 32'h1597cd39;
         473:    rdata = 32'h85930000;
         474:    rdata = 32'h85266265;
         475:    rdata = 32'h75a000ef;
         476:    rdata = 32'hc5314795;
         477:    rdata = 32'h00001597;
         478:    rdata = 32'h62058593;
         479:    rdata = 32'h00ef8526;
         480:    rdata = 32'h47997480;
         481:    rdata = 32'h1597cd0d;
         482:    rdata = 32'h85930000;
         483:    rdata = 32'h852661a5;
         484:    rdata = 32'h736000ef;
         485:    rdata = 32'hc505479d;
         486:    rdata = 32'h00001597;
         487:    rdata = 32'h61858593;
         488:    rdata = 32'h00ef8526;
         489:    rdata = 32'h47a17240;
         490:    rdata = 32'h1597c919;
         491:    rdata = 32'h85930000;
         492:    rdata = 32'h85266125;
         493:    rdata = 32'h712000ef;
         494:    rdata = 32'hc11147a5;
         495:    rdata = 32'hc01c47a9;
         496:    rdata = 32'h1101b7a9;
         497:    rdata = 32'hc84acc22;
         498:    rdata = 32'hc452c64e;
         499:    rdata = 32'hca26ce06;
         500:    rdata = 32'h8413892e;
         501:    rdata = 32'h498100c5;
         502:    rdata = 32'h27834a05;
         503:    rdata = 32'hd8630049;
         504:    rdata = 32'h049302f9;
         505:    rdata = 32'h85260184;
         506:    rdata = 32'h00ef0985;
         507:    rdata = 32'hc9090150;
         508:    rdata = 32'hff442e23;
         509:    rdata = 32'h00ef8526;
         510:    rdata = 32'hc00803f0;
         511:    rdata = 32'hbff18426;
         512:    rdata = 32'hfe042e23;
         513:    rdata = 32'h852285a6;
         514:    rdata = 32'h690000ef;
         515:    rdata = 32'h40f2bfc5;
         516:    rdata = 32'h44d24462;
         517:    rdata = 32'h49b24942;
         518:    rdata = 32'h61054a22;
         519:    rdata = 32'h11418082;
         520:    rdata = 32'hc422c606;
         521:    rdata = 32'hc04ac226;
         522:    rdata = 32'h84ae842a;
         523:    rdata = 32'h22238932;
         524:    rdata = 32'h06130005;
         525:    rdata = 32'h45810900;
         526:    rdata = 32'h00ef0521;
         527:    rdata = 32'h862273b0;
         528:    rdata = 32'h852685ca;
         529:    rdata = 32'h405c3591;
         530:    rdata = 32'h47adeb91;
         531:    rdata = 32'h40b2c01c;
         532:    rdata = 32'h44228522;
         533:    rdata = 32'h49024492;
         534:    rdata = 32'h80820141;
         535:    rdata = 32'h852685a2;
         536:    rdata = 32'h85a23561;
         537:    rdata = 32'h3fb18526;
         538:    rdata = 32'h7119b7dd;
         539:    rdata = 32'h006885aa;
         540:    rdata = 32'h251dde86;
         541:    rdata = 32'h00001597;
         542:    rdata = 32'h42058593;
         543:    rdata = 32'h25350068;
         544:    rdata = 32'hf517006c;
         545:    rdata = 32'h0513000e;
         546:    rdata = 32'h00ef7f65;
         547:    rdata = 32'h50f60a50;
         548:    rdata = 32'h80826109;
         549:    rdata = 32'h85aa1101;
         550:    rdata = 32'hce060048;
         551:    rdata = 32'h00482d5d;
         552:    rdata = 32'h40f237e9;
         553:    rdata = 32'h80826105;
         554:    rdata = 32'h85aa1101;
         555:    rdata = 32'hce060048;
         556:    rdata = 32'h708000ef;
         557:    rdata = 32'h3f550048;
         558:    rdata = 32'h610540f2;
         559:    rdata = 32'h71198082;
         560:    rdata = 32'h842edca2;
         561:    rdata = 32'h006885aa;
         562:    rdata = 32'h23f9de86;
         563:    rdata = 32'h00001597;
         564:    rdata = 32'h52458593;
         565:    rdata = 32'h2bd10068;
         566:    rdata = 32'h006885a2;
         567:    rdata = 32'h159723f9;
         568:    rdata = 32'h85930000;
         569:    rdata = 32'h00683b65;
         570:    rdata = 32'h006c23c9;
         571:    rdata = 32'h000ef517;
         572:    rdata = 32'h78c50513;
         573:    rdata = 32'h03b000ef;
         574:    rdata = 32'h546650f6;
         575:    rdata = 32'h80826109;
         576:    rdata = 32'hcc221101;
         577:    rdata = 32'h0048842a;
         578:    rdata = 32'h25a1ce06;
         579:    rdata = 32'h8522004c;
         580:    rdata = 32'h40f2377d;
         581:    rdata = 32'h61054462;
         582:    rdata = 32'h11018082;
         583:    rdata = 32'h842acc22;
         584:    rdata = 32'hce060048;
         585:    rdata = 32'h004c2d51;
         586:    rdata = 32'h3f518522;
         587:    rdata = 32'h446240f2;
         588:    rdata = 32'h80826105;
         589:    rdata = 32'hdaa67119;
         590:    rdata = 32'h85aa84ae;
         591:    rdata = 32'hde860068;
         592:    rdata = 32'h8432dca2;
         593:    rdata = 32'h15972b91;
         594:    rdata = 32'h85930000;
         595:    rdata = 32'h00684ae5;
         596:    rdata = 32'h85a62ba9;
         597:    rdata = 32'h2b910068;
         598:    rdata = 32'h00001597;
         599:    rdata = 32'h4a058593;
         600:    rdata = 32'h23a10068;
         601:    rdata = 32'h006885a2;
         602:    rdata = 32'h15972389;
         603:    rdata = 32'h85930000;
         604:    rdata = 32'h006832a5;
         605:    rdata = 32'h006c2b1d;
         606:    rdata = 32'h000ef517;
         607:    rdata = 32'h70050513;
         608:    rdata = 32'h7ae000ef;
         609:    rdata = 32'h546650f6;
         610:    rdata = 32'h610954d6;
         611:    rdata = 32'h71798082;
         612:    rdata = 32'h842ad422;
         613:    rdata = 32'hd6060028;
         614:    rdata = 32'h84b2d226;
         615:    rdata = 32'h85a62d31;
         616:    rdata = 32'h2b450848;
         617:    rdata = 32'h002c0850;
         618:    rdata = 32'h37698522;
         619:    rdata = 32'h542250b2;
         620:    rdata = 32'h61455492;
         621:    rdata = 32'h71798082;
         622:    rdata = 32'h842ad422;
         623:    rdata = 32'hd6060028;
         624:    rdata = 32'h84b2d226;
         625:    rdata = 32'h85a62bd5;
         626:    rdata = 32'h23fd0848;
         627:    rdata = 32'h002c0850;
         628:    rdata = 32'h378d8522;
         629:    rdata = 32'h542250b2;
         630:    rdata = 32'h61455492;
         631:    rdata = 32'h11018082;
         632:    rdata = 32'h842acc22;
         633:    rdata = 32'h000ef517;
         634:    rdata = 32'h65c50513;
         635:    rdata = 32'hca26ce06;
         636:    rdata = 32'hc64ec84a;
         637:    rdata = 32'h00efc452;
         638:    rdata = 32'hf51731b0;
         639:    rdata = 32'h0513000e;
         640:    rdata = 32'h00ef6465;
         641:    rdata = 32'hf4972310;
         642:    rdata = 32'h8493000e;
         643:    rdata = 32'h852663a4;
         644:    rdata = 32'h22f000ef;
         645:    rdata = 32'h44fddd6d;
         646:    rdata = 32'h000ef917;
         647:    rdata = 32'h62890913;
         648:    rdata = 32'h000efa17;
         649:    rdata = 32'h604a0a13;
         650:    rdata = 32'h854a59fd;
         651:    rdata = 32'h207000ef;
         652:    rdata = 32'h00ef854a;
         653:    rdata = 32'hdd6d20d0;
         654:    rdata = 32'h00649593;
         655:    rdata = 32'h855295a2;
         656:    rdata = 32'h00ef14fd;
         657:    rdata = 32'h92e31a10;
         658:    rdata = 32'h40f2ff34;
         659:    rdata = 32'h44628522;
         660:    rdata = 32'h494244d2;
         661:    rdata = 32'h4a2249b2;
         662:    rdata = 32'h80826105;
         663:    rdata = 32'hcc221101;
         664:    rdata = 32'hf517842a;
         665:    rdata = 32'h0513000e;
         666:    rdata = 32'hce065de5;
         667:    rdata = 32'h00efc62e;
         668:    rdata = 32'hf5172bd0;
         669:    rdata = 32'h0513000e;
         670:    rdata = 32'h00ef5ce5;
         671:    rdata = 32'h45b21b90;
         672:    rdata = 32'h3fb18522;
         673:    rdata = 32'h852240f2;
         674:    rdata = 32'h61054462;
         675:    rdata = 32'h715d8082;
         676:    rdata = 32'h872e878a;
         677:    rdata = 32'hc4a2c686;
         678:    rdata = 32'h85bec2a6;
         679:    rdata = 32'h00e79023;
         680:    rdata = 32'h07890094;
         681:    rdata = 32'hfed79ce3;
         682:    rdata = 32'h000ef517;
         683:    rdata = 32'h57c50513;
         684:    rdata = 32'h12b000ef;
         685:    rdata = 32'h000ef517;
         686:    rdata = 32'h58c50513;
         687:    rdata = 32'h255000ef;
         688:    rdata = 32'h000ef517;
         689:    rdata = 32'h58050513;
         690:    rdata = 32'h16b000ef;
         691:    rdata = 32'h000ef417;
         692:    rdata = 32'h57440413;
         693:    rdata = 32'h00ef8522;
         694:    rdata = 32'hdd6d1690;
         695:    rdata = 32'h02000413;
         696:    rdata = 32'h000ef497;
         697:    rdata = 32'h56048493;
         698:    rdata = 32'h00ef8526;
         699:    rdata = 32'h85261490;
         700:    rdata = 32'h14f000ef;
         701:    rdata = 32'h147ddd6d;
         702:    rdata = 32'h40b6f865;
         703:    rdata = 32'h44964426;
         704:    rdata = 32'h80826161;
         705:    rdata = 32'hc6061141;
         706:    rdata = 32'hf5173759;
         707:    rdata = 32'h0513000e;
         708:    rdata = 32'h00ef5365;
         709:    rdata = 32'h40b220d0;
         710:    rdata = 32'h000ef517;
         711:    rdata = 32'h52850513;
         712:    rdata = 32'h006f0141;
         713:    rdata = 32'h11011110;
         714:    rdata = 32'h000ef517;
         715:    rdata = 32'h51850513;
         716:    rdata = 32'hcc22ce06;
         717:    rdata = 32'hc84aca26;
         718:    rdata = 32'hc64e84ae;
         719:    rdata = 32'h1d5000ef;
         720:    rdata = 32'h000ef517;
         721:    rdata = 32'h50050513;
         722:    rdata = 32'h0eb000ef;
         723:    rdata = 32'h000ef417;
         724:    rdata = 32'h4f440413;
         725:    rdata = 32'h00ef8522;
         726:    rdata = 32'hdd6d0e90;
         727:    rdata = 32'h7c048413;
         728:    rdata = 32'h000ef997;
         729:    rdata = 32'h4c498993;
         730:    rdata = 32'h000ef917;
         731:    rdata = 32'h4d890913;
         732:    rdata = 32'h85a2854e;
         733:    rdata = 32'h067000ef;
         734:    rdata = 32'h00ef854a;
         735:    rdata = 32'h854a0b90;
         736:    rdata = 32'h0bf000ef;
         737:    rdata = 32'h0793dd6d;
         738:    rdata = 32'h9963fc04;
         739:    rdata = 32'h40f20084;
         740:    rdata = 32'h44d24462;
         741:    rdata = 32'h49b24942;
         742:    rdata = 32'h80826105;
         743:    rdata = 32'hbfc9843e;
         744:    rdata = 32'hc6061141;
         745:    rdata = 32'hf5173749;
         746:    rdata = 32'h0513000e;
         747:    rdata = 32'h00ef49a5;
         748:    rdata = 32'h40b21710;
         749:    rdata = 32'h000ef517;
         750:    rdata = 32'h48c50513;
         751:    rdata = 32'h006f0141;
         752:    rdata = 32'h71390750;
         753:    rdata = 32'hd452737d;
         754:    rdata = 32'h81030313;
         755:    rdata = 32'hdc226a09;
         756:    rdata = 32'hd84ada26;
         757:    rdata = 32'hd256d64e;
         758:    rdata = 32'hce5ed05a;
         759:    rdata = 32'hde06cc62;
         760:    rdata = 32'h800a0793;
         761:    rdata = 32'h978a911a;
         762:    rdata = 32'h84b3747d;
         763:    rdata = 32'h892a0087;
         764:    rdata = 32'h45816605;
         765:    rdata = 32'h00ef8526;
         766:    rdata = 32'h079337f0;
         767:    rdata = 32'h0413800a;
         768:    rdata = 32'h978a8004;
         769:    rdata = 32'h943e6a05;
         770:    rdata = 32'h880a0a13;
         771:    rdata = 32'h89934b01;
         772:    rdata = 32'h0b938004;
         773:    rdata = 32'h8aa60804;
         774:    rdata = 32'h0c139a22;
         775:    rdata = 32'h854a0800;
         776:    rdata = 32'h080b4433;
         777:    rdata = 32'h3df985a2;
         778:    rdata = 32'h85ca854e;
         779:    rdata = 32'h855e3d05;
         780:    rdata = 32'h0e138826;
         781:    rdata = 32'h0693f805;
         782:    rdata = 32'h03131808;
         783:    rdata = 32'h07130405;
         784:    rdata = 32'h07931008;
         785:    rdata = 32'h05930808;
         786:    rdata = 32'h88aafc05;
         787:    rdata = 32'h5e838642;
         788:    rdata = 32'h5f03000e;
         789:    rdata = 32'h76630026;
         790:    rdata = 32'h102301df;
         791:    rdata = 32'h11230086;
         792:    rdata = 32'h5e8301d6;
         793:    rdata = 32'h5f03002e;
         794:    rdata = 32'h76630066;
         795:    rdata = 32'h122301df;
         796:    rdata = 32'h13230086;
         797:    rdata = 32'h5e8301d6;
         798:    rdata = 32'h5f03004e;
         799:    rdata = 32'h766300a6;
         800:    rdata = 32'h142301df;
         801:    rdata = 32'h15230086;
         802:    rdata = 32'h5e8301d6;
         803:    rdata = 32'h5f03006e;
         804:    rdata = 32'h766300e6;
         805:    rdata = 32'h162301df;
         806:    rdata = 32'h17230086;
         807:    rdata = 32'hde8301d6;
         808:    rdata = 32'hdf030005;
         809:    rdata = 32'h76630027;
         810:    rdata = 32'h902301df;
         811:    rdata = 32'h91230087;
         812:    rdata = 32'hde8301d7;
         813:    rdata = 32'hdf030025;
         814:    rdata = 32'h76630067;
         815:    rdata = 32'h922301df;
         816:    rdata = 32'h93230087;
         817:    rdata = 32'hde8301d7;
         818:    rdata = 32'hdf030045;
         819:    rdata = 32'h766300a7;
         820:    rdata = 32'h942301df;
         821:    rdata = 32'h95230087;
         822:    rdata = 32'hde8301d7;
         823:    rdata = 32'hdf030065;
         824:    rdata = 32'h766300e7;
         825:    rdata = 32'h962301df;
         826:    rdata = 32'h97230087;
         827:    rdata = 32'hde8301d7;
         828:    rdata = 32'h5f030008;
         829:    rdata = 32'h76630027;
         830:    rdata = 32'h102301df;
         831:    rdata = 32'h11230087;
         832:    rdata = 32'hde8301d7;
         833:    rdata = 32'h5f030028;
         834:    rdata = 32'h76630067;
         835:    rdata = 32'h122301df;
         836:    rdata = 32'h13230087;
         837:    rdata = 32'hde8301d7;
         838:    rdata = 32'h5f030048;
         839:    rdata = 32'h766300a7;
         840:    rdata = 32'h142301df;
         841:    rdata = 32'h15230087;
         842:    rdata = 32'hde8301d7;
         843:    rdata = 32'h5f030068;
         844:    rdata = 32'h766300e7;
         845:    rdata = 32'h162301df;
         846:    rdata = 32'h17230087;
         847:    rdata = 32'h5e8301d7;
         848:    rdata = 32'hdf030003;
         849:    rdata = 32'h76630026;
         850:    rdata = 32'h902301df;
         851:    rdata = 32'h91230086;
         852:    rdata = 32'h5e8301d6;
         853:    rdata = 32'hdf030023;
         854:    rdata = 32'h76630066;
         855:    rdata = 32'h922301df;
         856:    rdata = 32'h93230086;
         857:    rdata = 32'h5e8301d6;
         858:    rdata = 32'hdf030043;
         859:    rdata = 32'h766300a6;
         860:    rdata = 32'h942301df;
         861:    rdata = 32'h95230086;
         862:    rdata = 32'h5e8301d6;
         863:    rdata = 32'hdf030063;
         864:    rdata = 32'h766300e6;
         865:    rdata = 32'h962301df;
         866:    rdata = 32'h97230086;
         867:    rdata = 32'h05a101d6;
         868:    rdata = 32'h06410e21;
         869:    rdata = 32'h032106c1;
         870:    rdata = 32'h08a10741;
         871:    rdata = 32'h98e307c1;
         872:    rdata = 32'h8513eaa5;
         873:    rdata = 32'h08131005;
         874:    rdata = 32'h14e32008;
         875:    rdata = 32'h0b05e945;
         876:    rdata = 32'he78b17e3;
         877:    rdata = 32'h777d6789;
         878:    rdata = 32'h80078793;
         879:    rdata = 32'h0713978a;
         880:    rdata = 32'h973e8007;
         881:    rdata = 32'h94be6785;
         882:    rdata = 32'h86ba87d6;
         883:    rdata = 32'h080a8a93;
         884:    rdata = 32'h0007d603;
         885:    rdata = 32'h06890791;
         886:    rdata = 32'hfec69f23;
         887:    rdata = 32'hfefa9ae3;
         888:    rdata = 32'h04070713;
         889:    rdata = 32'hfe9a92e3;
         890:    rdata = 32'h75fd6789;
         891:    rdata = 32'h80078793;
         892:    rdata = 32'h8593978a;
         893:    rdata = 32'h854a8005;
         894:    rdata = 32'h335d95be;
         895:    rdata = 32'h03136305;
         896:    rdata = 32'h911a7f03;
         897:    rdata = 32'h546250f2;
         898:    rdata = 32'h594254d2;
         899:    rdata = 32'h5a2259b2;
         900:    rdata = 32'h5b025a92;
         901:    rdata = 32'h4c624bf2;
         902:    rdata = 32'h80826121;
         903:    rdata = 32'h03000713;
         904:    rdata = 32'h00054783;
         905:    rdata = 32'h00e79463;
         906:    rdata = 32'hbfdd0505;
         907:    rdata = 32'h157de391;
         908:    rdata = 32'h47038082;
         909:    rdata = 32'h07930005;
         910:    rdata = 32'h136302d0;
         911:    rdata = 32'h050500f7;
         912:    rdata = 32'h47834725;
         913:    rdata = 32'h87930005;
         914:    rdata = 32'hf793fd07;
         915:    rdata = 32'h68630ff7;
         916:    rdata = 32'h478300f7;
         917:    rdata = 32'h05050015;
         918:    rdata = 32'h4505f7ed;
         919:    rdata = 32'h45018082;
         920:    rdata = 32'h05098082;
         921:    rdata = 32'h461546a5;
         922:    rdata = 32'h00054783;
         923:    rdata = 32'hfd078713;
         924:    rdata = 32'h0ff77713;
         925:    rdata = 32'h00e6fa63;
         926:    rdata = 32'hfdf7f793;
         927:    rdata = 32'hfbf78793;
         928:    rdata = 32'h0ff7f793;
         929:    rdata = 32'h00f66863;
         930:    rdata = 32'h00154783;
         931:    rdata = 32'hffe90505;
         932:    rdata = 32'h80824505;
         933:    rdata = 32'h80824501;
         934:    rdata = 32'hc70387aa;
         935:    rdata = 32'h05850005;
         936:    rdata = 32'h8fa30785;
         937:    rdata = 32'hfb75fee7;
         938:    rdata = 32'h87aa8082;
         939:    rdata = 32'h0007c683;
         940:    rdata = 32'h0785873e;
         941:    rdata = 32'hc783fee5;
         942:    rdata = 32'h05850005;
         943:    rdata = 32'h0fa30705;
         944:    rdata = 32'hfbf5fef7;
         945:    rdata = 32'h47838082;
         946:    rdata = 32'hc7030005;
         947:    rdata = 32'h87630005;
         948:    rdata = 32'h557d00e7;
         949:    rdata = 32'h00e7e963;
         950:    rdata = 32'h80824505;
         951:    rdata = 32'h0505c781;
         952:    rdata = 32'hb7d50585;
         953:    rdata = 32'h80824501;
         954:    rdata = 32'h450187aa;
         955:    rdata = 32'h00a78733;
         956:    rdata = 32'h00074703;
         957:    rdata = 32'h0505c319;
         958:    rdata = 32'h8082bfd5;
         959:    rdata = 32'h0c634789;
         960:    rdata = 32'h479102f6;
         961:    rdata = 32'h02f60d63;
         962:    rdata = 32'h47814705;
         963:    rdata = 32'h00e61463;
         964:    rdata = 32'h06400793;
         965:    rdata = 32'hcb8d4629;
         966:    rdata = 32'h02f5d733;
         967:    rdata = 32'h76930505;
         968:    rdata = 32'h86b30ff7;
         969:    rdata = 32'h071302f6;
         970:    rdata = 32'h0fa30307;
         971:    rdata = 32'hd7b3fee5;
         972:    rdata = 32'h8d9502c7;
         973:    rdata = 32'h6789b7cd;
         974:    rdata = 32'h71078793;
         975:    rdata = 32'hd7b7bfe1;
         976:    rdata = 32'h87933b9a;
         977:    rdata = 32'hb7f9a007;
         978:    rdata = 32'h00050023;
         979:    rdata = 32'h46058082;
         980:    rdata = 32'h1101b775;
         981:    rdata = 32'h4611cc22;
         982:    rdata = 32'h0048842a;
         983:    rdata = 32'h3f79ce06;
         984:    rdata = 32'h3d6d0048;
         985:    rdata = 32'h852285aa;
         986:    rdata = 32'h40f23f05;
         987:    rdata = 32'h61054462;
         988:    rdata = 32'h07938082;
         989:    rdata = 32'h06060300;
         990:    rdata = 32'h0ff67613;
         991:    rdata = 32'h00f50023;
         992:    rdata = 32'h07800793;
         993:    rdata = 32'h00f500a3;
         994:    rdata = 32'h87b24825;
         995:    rdata = 32'hf713c385;
         996:    rdata = 32'h069300f5;
         997:    rdata = 32'h64630577;
         998:    rdata = 32'h069300e8;
         999:    rdata = 32'h07330307;
        1000:    rdata = 32'h00a300f5;
        1001:    rdata = 32'h819100d7;
        1002:    rdata = 32'hb7cd17fd;
        1003:    rdata = 32'h01239532;
        1004:    rdata = 32'h80820005;
        1005:    rdata = 32'hbf754605;
        1006:    rdata = 32'hbf654611;
        1007:    rdata = 32'hcc221101;
        1008:    rdata = 32'h842ace06;
        1009:    rdata = 32'h0205d563;
        1010:    rdata = 32'h02d00713;
        1011:    rdata = 32'h00e50023;
        1012:    rdata = 32'h40b005b3;
        1013:    rdata = 32'h00484611;
        1014:    rdata = 32'h00483715;
        1015:    rdata = 32'h85aa3581;
        1016:    rdata = 32'h00140513;
        1017:    rdata = 32'h40f23d55;
        1018:    rdata = 32'h61054462;
        1019:    rdata = 32'h46118082;
        1020:    rdata = 32'h37290048;
        1021:    rdata = 32'h351d0048;
        1022:    rdata = 32'h852285aa;
        1023:    rdata = 32'h1141b7e5;
        1024:    rdata = 32'hc606c422;
        1025:    rdata = 32'h3535842a;
        1026:    rdata = 32'h4703e115;
        1027:    rdata = 32'h07930004;
        1028:    rdata = 32'h1d630300;
        1029:    rdata = 32'h470300f7;
        1030:    rdata = 32'h07930014;
        1031:    rdata = 32'h17630780;
        1032:    rdata = 32'h852200f7;
        1033:    rdata = 32'h40b24422;
        1034:    rdata = 32'hbd250141;
        1035:    rdata = 32'h442240b2;
        1036:    rdata = 32'h80820141;
        1037:    rdata = 32'hc4221141;
        1038:    rdata = 32'h842ac606;
        1039:    rdata = 32'h47833bdd;
        1040:    rdata = 32'hc91d0004;
        1041:    rdata = 32'h02d00693;
        1042:    rdata = 32'h94634701;
        1043:    rdata = 32'h872a00d7;
        1044:    rdata = 32'h45010405;
        1045:    rdata = 32'h46834629;
        1046:    rdata = 32'hca810004;
        1047:    rdata = 32'h02c507b3;
        1048:    rdata = 32'hfd068513;
        1049:    rdata = 32'h953e0405;
        1050:    rdata = 32'hc319b7fd;
        1051:    rdata = 32'h40a00533;
        1052:    rdata = 32'h442240b2;
        1053:    rdata = 32'h80820141;
        1054:    rdata = 32'h03000713;
        1055:    rdata = 32'h04e79663;
        1056:    rdata = 32'h00144703;
        1057:    rdata = 32'h07800793;
        1058:    rdata = 32'h04f71063;
        1059:    rdata = 32'h3bd18522;
        1060:    rdata = 32'h0409cd05;
        1061:    rdata = 32'h07134501;
        1062:    rdata = 32'h06930600;
        1063:    rdata = 32'h47830400;
        1064:    rdata = 32'hd7f90004;
        1065:    rdata = 32'h00f77a63;
        1066:    rdata = 32'hfa978793;
        1067:    rdata = 32'h0ff7f793;
        1068:    rdata = 32'h8d5d0512;
        1069:    rdata = 32'hb7e50405;
        1070:    rdata = 32'h00f6f563;
        1071:    rdata = 32'hfc978793;
        1072:    rdata = 32'h8793b7f5;
        1073:    rdata = 32'hb7ddfd07;
        1074:    rdata = 32'hdeadc537;
        1075:    rdata = 32'heef50513;
        1076:    rdata = 32'h7793b745;
        1077:    rdata = 32'h8793fdf5;
        1078:    rdata = 32'hf793fbf7;
        1079:    rdata = 32'h47650ff7;
        1080:    rdata = 32'h00f77763;
        1081:    rdata = 32'hfd050513;
        1082:    rdata = 32'h00a53513;
        1083:    rdata = 32'h45058082;
        1084:    rdata = 32'h11418082;
        1085:    rdata = 32'h0613c422;
        1086:    rdata = 32'h842a0640;
        1087:    rdata = 32'h000ef517;
        1088:    rdata = 32'hf6450513;
        1089:    rdata = 32'h214dc606;
        1090:    rdata = 32'h852240b2;
        1091:    rdata = 32'h01414422;
        1092:    rdata = 32'h11418082;
        1093:    rdata = 32'h842ac422;
        1094:    rdata = 32'h000ef517;
        1095:    rdata = 32'hf4850513;
        1096:    rdata = 32'h29e5c606;
        1097:    rdata = 32'h852240b2;
        1098:    rdata = 32'h01414422;
        1099:    rdata = 32'h11418082;
        1100:    rdata = 32'h842ac422;
        1101:    rdata = 32'h000ef517;
        1102:    rdata = 32'hf2c50513;
        1103:    rdata = 32'h29f1c606;
        1104:    rdata = 32'h852240b2;
        1105:    rdata = 32'h01414422;
        1106:    rdata = 32'h418c8082;
        1107:    rdata = 32'hcc221101;
        1108:    rdata = 32'h0048842a;
        1109:    rdata = 32'h359dce06;
        1110:    rdata = 32'hf517004c;
        1111:    rdata = 32'h0513000e;
        1112:    rdata = 32'h2965f065;
        1113:    rdata = 32'h852240f2;
        1114:    rdata = 32'h61054462;
        1115:    rdata = 32'h71758082;
        1116:    rdata = 32'hc326c522;
        1117:    rdata = 32'hdecec14a;
        1118:    rdata = 32'hc706dcd2;
        1119:    rdata = 32'h892e84aa;
        1120:    rdata = 32'h000ef417;
        1121:    rdata = 32'hee040413;
        1122:    rdata = 32'h00001a17;
        1123:    rdata = 32'hc68a0a13;
        1124:    rdata = 32'h00001997;
        1125:    rdata = 32'hc6c98993;
        1126:    rdata = 32'h852285ca;
        1127:    rdata = 32'h85d229bd;
        1128:    rdata = 32'h29a58522;
        1129:    rdata = 32'h8526006c;
        1130:    rdata = 32'h006837a9;
        1131:    rdata = 32'he5093d89;
        1132:    rdata = 32'h852285ce;
        1133:    rdata = 32'hb7cd219d;
        1134:    rdata = 32'h3dad0068;
        1135:    rdata = 32'h442a40ba;
        1136:    rdata = 32'h490a449a;
        1137:    rdata = 32'h5a6659f6;
        1138:    rdata = 32'h80826149;
        1139:    rdata = 32'hb0002573;
        1140:    rdata = 32'hb80025f3;
        1141:    rdata = 32'h00018082;
        1142:    rdata = 32'h00010001;
        1143:    rdata = 32'h00010001;
        1144:    rdata = 32'h15fd0001;
        1145:    rdata = 32'h8082f9ed;
        1146:    rdata = 32'h300462f3;
        1147:    rdata = 32'h72f38082;
        1148:    rdata = 32'h80823004;
        1149:    rdata = 32'h62c1c10c;
        1150:    rdata = 32'h3042a2f3;
        1151:    rdata = 32'h20238082;
        1152:    rdata = 32'h62c10005;
        1153:    rdata = 32'h3042b2f3;
        1154:    rdata = 32'hc14c8082;
        1155:    rdata = 32'h000202b7;
        1156:    rdata = 32'h3042a2f3;
        1157:    rdata = 32'h22238082;
        1158:    rdata = 32'h02b70005;
        1159:    rdata = 32'hb2f30002;
        1160:    rdata = 32'h80823042;
        1161:    rdata = 32'hcc3e7139;
        1162:    rdata = 32'hdc16de06;
        1163:    rdata = 32'hd81eda1a;
        1164:    rdata = 32'hd42ed62a;
        1165:    rdata = 32'hd036d232;
        1166:    rdata = 32'hca42ce3a;
        1167:    rdata = 32'hc672c846;
        1168:    rdata = 32'hc27ac476;
        1169:    rdata = 32'hf797c07e;
        1170:    rdata = 32'ha783000e;
        1171:    rdata = 32'h9782e367;
        1172:    rdata = 32'h52e250f2;
        1173:    rdata = 32'h53c25352;
        1174:    rdata = 32'h55a25532;
        1175:    rdata = 32'h56825612;
        1176:    rdata = 32'h47e24772;
        1177:    rdata = 32'h48c24852;
        1178:    rdata = 32'h4ea24e32;
        1179:    rdata = 32'h4f824f12;
        1180:    rdata = 32'h00736121;
        1181:    rdata = 32'h71393020;
        1182:    rdata = 32'hde06cc3e;
        1183:    rdata = 32'hda1adc16;
        1184:    rdata = 32'hd62ad81e;
        1185:    rdata = 32'hd232d42e;
        1186:    rdata = 32'hce3ad036;
        1187:    rdata = 32'hc846ca42;
        1188:    rdata = 32'hc476c672;
        1189:    rdata = 32'hc07ec27a;
        1190:    rdata = 32'h000ef797;
        1191:    rdata = 32'hde87a783;
        1192:    rdata = 32'h50f29782;
        1193:    rdata = 32'h535252e2;
        1194:    rdata = 32'h553253c2;
        1195:    rdata = 32'h561255a2;
        1196:    rdata = 32'h47725682;
        1197:    rdata = 32'h485247e2;
        1198:    rdata = 32'h4e3248c2;
        1199:    rdata = 32'h4f124ea2;
        1200:    rdata = 32'h61214f82;
        1201:    rdata = 32'h30200073;
        1202:    rdata = 32'h00458793;
        1203:    rdata = 32'h8793c15c;
        1204:    rdata = 32'hc51c0085;
        1205:    rdata = 32'h00c58793;
        1206:    rdata = 32'h8793c55c;
        1207:    rdata = 32'hc91c0105;
        1208:    rdata = 32'h01458793;
        1209:    rdata = 32'h8793c95c;
        1210:    rdata = 32'hc10c0185;
        1211:    rdata = 32'h8793cd1c;
        1212:    rdata = 32'h859301c5;
        1213:    rdata = 32'hcd5c0205;
        1214:    rdata = 32'h8082d10c;
        1215:    rdata = 32'h8a05511c;
        1216:    rdata = 32'h00b61633;
        1217:    rdata = 32'h97b3439c;
        1218:    rdata = 32'h8e5d48b7;
        1219:    rdata = 32'hc390511c;
        1220:    rdata = 32'h511c8082;
        1221:    rdata = 32'h47854388;
        1222:    rdata = 32'h00b797b3;
        1223:    rdata = 32'h35338d7d;
        1224:    rdata = 32'h808200a0;
        1225:    rdata = 32'h4388455c;
        1226:    rdata = 32'h97b34785;
        1227:    rdata = 32'h8d7d00b7;
        1228:    rdata = 32'h00a03533;
        1229:    rdata = 32'h451c8082;
        1230:    rdata = 32'h8e3d439c;
        1231:    rdata = 32'h8e3d8e6d;
        1232:    rdata = 32'hc390451c;
        1233:    rdata = 32'h47858082;
        1234:    rdata = 32'h00b61633;
        1235:    rdata = 32'h00b795b3;
        1236:    rdata = 32'h1141b7dd;
        1237:    rdata = 32'hc226c422;
        1238:    rdata = 32'h842ac606;
        1239:    rdata = 32'h37d984ae;
        1240:    rdata = 32'h00154613;
        1241:    rdata = 32'h44228522;
        1242:    rdata = 32'h85a640b2;
        1243:    rdata = 32'h76134492;
        1244:    rdata = 32'h01410ff6;
        1245:    rdata = 32'h455cbfc9;
        1246:    rdata = 32'h55134388;
        1247:    rdata = 32'h80824915;
        1248:    rdata = 32'h4388455c;
        1249:    rdata = 32'h49055513;
        1250:    rdata = 32'h11418082;
        1251:    rdata = 32'h4601c226;
        1252:    rdata = 32'h45bd84ae;
        1253:    rdata = 32'hc606c422;
        1254:    rdata = 32'h378d842a;
        1255:    rdata = 32'h44228522;
        1256:    rdata = 32'h862640b2;
        1257:    rdata = 32'h45bd4492;
        1258:    rdata = 32'hbf710141;
        1259:    rdata = 32'h00858713;
        1260:    rdata = 32'h05058793;
        1261:    rdata = 32'hc91cc518;
        1262:    rdata = 32'h01058713;
        1263:    rdata = 32'h010107b7;
        1264:    rdata = 32'h8613c558;
        1265:    rdata = 32'h87130045;
        1266:    rdata = 32'h87931007;
        1267:    rdata = 32'hc10c2007;
        1268:    rdata = 32'hc958c150;
        1269:    rdata = 32'h0571cd1c;
        1270:    rdata = 32'h4548a81d;
        1271:    rdata = 32'h04000613;
        1272:    rdata = 32'h87aaaca5;
        1273:    rdata = 32'h4b8c852e;
        1274:    rdata = 32'h04000613;
        1275:    rdata = 32'h495ca4b5;
        1276:    rdata = 32'hc3984198;
        1277:    rdata = 32'h41d8495c;
        1278:    rdata = 32'h4598c3d8;
        1279:    rdata = 32'hc798495c;
        1280:    rdata = 32'h495c45d8;
        1281:    rdata = 32'h8082c7d8;
        1282:    rdata = 32'hc38c4d1c;
        1283:    rdata = 32'hc10c8082;
        1284:    rdata = 32'h15b7c150;
        1285:    rdata = 32'h06130101;
        1286:    rdata = 32'h05214000;
        1287:    rdata = 32'h4118a42d;
        1288:    rdata = 32'h0015c593;
        1289:    rdata = 32'h0015f793;
        1290:    rdata = 32'h99f9430c;
        1291:    rdata = 32'hc30c8ddd;
        1292:    rdata = 32'h41188082;
        1293:    rdata = 32'he793431c;
        1294:    rdata = 32'hc31c0027;
        1295:    rdata = 32'h415c8082;
        1296:    rdata = 32'h89054388;
        1297:    rdata = 32'h71398082;
        1298:    rdata = 32'h4411dc22;
        1299:    rdata = 32'h02864433;
        1300:    rdata = 32'hda264118;
        1301:    rdata = 32'hd64ed84a;
        1302:    rdata = 32'hd256d452;
        1303:    rdata = 32'hcc62ce5e;
        1304:    rdata = 32'hd05ade06;
        1305:    rdata = 32'h84aa431c;
        1306:    rdata = 32'h9bf989ae;
        1307:    rdata = 32'hc31c8932;
        1308:    rdata = 32'h4a814a01;
        1309:    rdata = 32'h0b934c11;
        1310:    rdata = 32'hd9630085;
        1311:    rdata = 32'h4781028a;
        1312:    rdata = 32'h01498633;
        1313:    rdata = 32'h00f606b3;
        1314:    rdata = 32'h0006c683;
        1315:    rdata = 32'h973e0078;
        1316:    rdata = 32'h00d70023;
        1317:    rdata = 32'h97e30785;
        1318:    rdata = 32'h4b32ff87;
        1319:    rdata = 32'h855e85d2;
        1320:    rdata = 32'h20232275;
        1321:    rdata = 32'h0a850165;
        1322:    rdata = 32'hbfc10a11;
        1323:    rdata = 32'h54334581;
        1324:    rdata = 32'h15930ab4;
        1325:    rdata = 32'h05330024;
        1326:    rdata = 32'h0a6340b9;
        1327:    rdata = 32'h478102b9;
        1328:    rdata = 32'h4701468d;
        1329:    rdata = 32'h00a7d763;
        1330:    rdata = 32'h00f58733;
        1331:    rdata = 32'h4703974e;
        1332:    rdata = 32'h00700007;
        1333:    rdata = 32'h0023963e;
        1334:    rdata = 32'h078500e6;
        1335:    rdata = 32'hfed793e3;
        1336:    rdata = 32'h000107a3;
        1337:    rdata = 32'h85134432;
        1338:    rdata = 32'h228d0084;
        1339:    rdata = 32'h4098c100;
        1340:    rdata = 32'he793431c;
        1341:    rdata = 32'hc31c0017;
        1342:    rdata = 32'h546250f2;
        1343:    rdata = 32'h594254d2;
        1344:    rdata = 32'h5a2259b2;
        1345:    rdata = 32'h5b025a92;
        1346:    rdata = 32'h4c624bf2;
        1347:    rdata = 32'h80826121;
        1348:    rdata = 32'h06700613;
        1349:    rdata = 32'h00000597;
        1350:    rdata = 32'h41458593;
        1351:    rdata = 32'h4625b72d;
        1352:    rdata = 32'h00000597;
        1353:    rdata = 32'h47058593;
        1354:    rdata = 32'h4625bf39;
        1355:    rdata = 32'h00000597;
        1356:    rdata = 32'h47058593;
        1357:    rdata = 32'h8793bf09;
        1358:    rdata = 32'hc10c0045;
        1359:    rdata = 32'h8793c15c;
        1360:    rdata = 32'h05b10085;
        1361:    rdata = 32'hc54cc51c;
        1362:    rdata = 32'h41188082;
        1363:    rdata = 32'he793431c;
        1364:    rdata = 32'hc31c0017;
        1365:    rdata = 32'h41188082;
        1366:    rdata = 32'h9bf9431c;
        1367:    rdata = 32'h8082c31c;
        1368:    rdata = 32'h431c4158;
        1369:    rdata = 32'hc31c9bf9;
        1370:    rdata = 32'h87938082;
        1371:    rdata = 32'hc15c0045;
        1372:    rdata = 32'h00858793;
        1373:    rdata = 32'h8793c51c;
        1374:    rdata = 32'hc55c00c5;
        1375:    rdata = 32'h01058793;
        1376:    rdata = 32'h47b1c91c;
        1377:    rdata = 32'h8823c10c;
        1378:    rdata = 32'h419c00f5;
        1379:    rdata = 32'h0017e793;
        1380:    rdata = 32'h8082c19c;
        1381:    rdata = 32'h439c415c;
        1382:    rdata = 32'hdfed8b85;
        1383:    rdata = 32'hc503455c;
        1384:    rdata = 32'h75130007;
        1385:    rdata = 32'h80820ff5;
        1386:    rdata = 32'hcc221101;
        1387:    rdata = 32'hc84aca26;
        1388:    rdata = 32'hc256c64e;
        1389:    rdata = 32'hce06c05a;
        1390:    rdata = 32'h84aac452;
        1391:    rdata = 32'h89b2892e;
        1392:    rdata = 32'h4aa94401;
        1393:    rdata = 32'h5f634b21;
        1394:    rdata = 32'h85260334;
        1395:    rdata = 32'h00890a33;
        1396:    rdata = 32'h002337d1;
        1397:    rdata = 32'h1f6300aa;
        1398:    rdata = 32'h00230155;
        1399:    rdata = 32'h4501000a;
        1400:    rdata = 32'h446240f2;
        1401:    rdata = 32'h494244d2;
        1402:    rdata = 32'h4a2249b2;
        1403:    rdata = 32'h4b024a92;
        1404:    rdata = 32'h80826105;
        1405:    rdata = 32'h01651463;
        1406:    rdata = 32'h1479c401;
        1407:    rdata = 32'hb7e10405;
        1408:    rdata = 32'hbfed547d;
        1409:    rdata = 32'hbfe94505;
        1410:    rdata = 32'h8023451c;
        1411:    rdata = 32'h415c00b7;
        1412:    rdata = 32'hd793439c;
        1413:    rdata = 32'hffe54817;
        1414:    rdata = 32'h11418082;
        1415:    rdata = 32'hc226c422;
        1416:    rdata = 32'h84aac606;
        1417:    rdata = 32'h4583842e;
        1418:    rdata = 32'hc5890004;
        1419:    rdata = 32'h04058526;
        1420:    rdata = 32'hbfd53fe1;
        1421:    rdata = 32'h442240b2;
        1422:    rdata = 32'h01414492;
        1423:    rdata = 32'h415c8082;
        1424:    rdata = 32'h89054388;
        1425:    rdata = 32'hc10c8082;
        1426:    rdata = 32'h8082c150;
        1427:    rdata = 32'h99f14108;
        1428:    rdata = 32'h8082952e;
        1429:    rdata = 32'h80824148;
        1430:    rdata = 32'h00a5c7b3;
        1431:    rdata = 32'h0037f793;
        1432:    rdata = 32'h00c508b3;
        1433:    rdata = 32'h06079263;
        1434:    rdata = 32'h00300793;
        1435:    rdata = 32'h04c7fe63;
        1436:    rdata = 32'h00357793;
        1437:    rdata = 32'h00050713;
        1438:    rdata = 32'h06079863;
        1439:    rdata = 32'hffc8f613;
        1440:    rdata = 32'hfe060793;
        1441:    rdata = 32'h08f76c63;
        1442:    rdata = 32'h02c77c63;
        1443:    rdata = 32'h00058693;
        1444:    rdata = 32'h00070793;
        1445:    rdata = 32'h0006a803;
        1446:    rdata = 32'h00478793;
        1447:    rdata = 32'h00468693;
        1448:    rdata = 32'hff07ae23;
        1449:    rdata = 32'hfec7e8e3;
        1450:    rdata = 32'hfff60793;
        1451:    rdata = 32'h40e787b3;
        1452:    rdata = 32'hffc7f793;
        1453:    rdata = 32'h00478793;
        1454:    rdata = 32'h00f70733;
        1455:    rdata = 32'h00f585b3;
        1456:    rdata = 32'h01176863;
        1457:    rdata = 32'h00008067;
        1458:    rdata = 32'h00050713;
        1459:    rdata = 32'hff157ce3;
        1460:    rdata = 32'h0005c783;
        1461:    rdata = 32'h00170713;
        1462:    rdata = 32'h00158593;
        1463:    rdata = 32'hfef70fa3;
        1464:    rdata = 32'hff1768e3;
        1465:    rdata = 32'h00008067;
        1466:    rdata = 32'h0005c683;
        1467:    rdata = 32'h00170713;
        1468:    rdata = 32'h00377793;
        1469:    rdata = 32'hfed70fa3;
        1470:    rdata = 32'h00158593;
        1471:    rdata = 32'hf80780e3;
        1472:    rdata = 32'h0005c683;
        1473:    rdata = 32'h00170713;
        1474:    rdata = 32'h00377793;
        1475:    rdata = 32'hfed70fa3;
        1476:    rdata = 32'h00158593;
        1477:    rdata = 32'hfc079ae3;
        1478:    rdata = 32'hf65ff06f;
        1479:    rdata = 32'h0045a683;
        1480:    rdata = 32'h0005a283;
        1481:    rdata = 32'h0085af83;
        1482:    rdata = 32'h00c5af03;
        1483:    rdata = 32'h0105ae83;
        1484:    rdata = 32'h0145ae03;
        1485:    rdata = 32'h0185a303;
        1486:    rdata = 32'h01c5a803;
        1487:    rdata = 32'h00d72223;
        1488:    rdata = 32'h0205a683;
        1489:    rdata = 32'h00572023;
        1490:    rdata = 32'h01f72423;
        1491:    rdata = 32'h01e72623;
        1492:    rdata = 32'h01d72823;
        1493:    rdata = 32'h01c72a23;
        1494:    rdata = 32'h00672c23;
        1495:    rdata = 32'h01072e23;
        1496:    rdata = 32'h02d72023;
        1497:    rdata = 32'h02470713;
        1498:    rdata = 32'h02458593;
        1499:    rdata = 32'hfaf768e3;
        1500:    rdata = 32'hf19ff06f;
        1501:    rdata = 32'h00f00313;
        1502:    rdata = 32'h00050713;
        1503:    rdata = 32'h02c37e63;
        1504:    rdata = 32'h00f77793;
        1505:    rdata = 32'h0a079063;
        1506:    rdata = 32'h08059263;
        1507:    rdata = 32'hff067693;
        1508:    rdata = 32'h00f67613;
        1509:    rdata = 32'h00e686b3;
        1510:    rdata = 32'h00b72023;
        1511:    rdata = 32'h00b72223;
        1512:    rdata = 32'h00b72423;
        1513:    rdata = 32'h00b72623;
        1514:    rdata = 32'h01070713;
        1515:    rdata = 32'hfed766e3;
        1516:    rdata = 32'h00061463;
        1517:    rdata = 32'h00008067;
        1518:    rdata = 32'h40c306b3;
        1519:    rdata = 32'h00269693;
        1520:    rdata = 32'h00000297;
        1521:    rdata = 32'h005686b3;
        1522:    rdata = 32'h00c68067;
        1523:    rdata = 32'h00b70723;
        1524:    rdata = 32'h00b706a3;
        1525:    rdata = 32'h00b70623;
        1526:    rdata = 32'h00b705a3;
        1527:    rdata = 32'h00b70523;
        1528:    rdata = 32'h00b704a3;
        1529:    rdata = 32'h00b70423;
        1530:    rdata = 32'h00b703a3;
        1531:    rdata = 32'h00b70323;
        1532:    rdata = 32'h00b702a3;
        1533:    rdata = 32'h00b70223;
        1534:    rdata = 32'h00b701a3;
        1535:    rdata = 32'h00b70123;
        1536:    rdata = 32'h00b700a3;
        1537:    rdata = 32'h00b70023;
        1538:    rdata = 32'h00008067;
        1539:    rdata = 32'h0ff5f593;
        1540:    rdata = 32'h00859693;
        1541:    rdata = 32'h00d5e5b3;
        1542:    rdata = 32'h01059693;
        1543:    rdata = 32'h00d5e5b3;
        1544:    rdata = 32'hf6dff06f;
        1545:    rdata = 32'h00279693;
        1546:    rdata = 32'h00000297;
        1547:    rdata = 32'h005686b3;
        1548:    rdata = 32'h00008293;
        1549:    rdata = 32'hfa0680e7;
        1550:    rdata = 32'h00028093;
        1551:    rdata = 32'hff078793;
        1552:    rdata = 32'h40f70733;
        1553:    rdata = 32'h00f60633;
        1554:    rdata = 32'hf6c378e3;
        1555:    rdata = 32'hf3dff06f;
        1556:    rdata = 32'h05971101;
        1557:    rdata = 32'h85930000;
        1558:    rdata = 32'hf51757e5;
        1559:    rdata = 32'h0513000e;
        1560:    rdata = 32'hce0681e5;
        1561:    rdata = 32'h8cbff0ef;
        1562:    rdata = 32'he0ef0068;
        1563:    rdata = 32'h40f2cfbf;
        1564:    rdata = 32'h61054501;
        1565:    rdata = 32'h05b78082;
        1566:    rdata = 32'he5170100;
        1567:    rdata = 32'h0513000e;
        1568:    rdata = 32'hf06f7865;
        1569:    rdata = 32'h05b7a47f;
        1570:    rdata = 32'he5170101;
        1571:    rdata = 32'h0513000e;
        1572:    rdata = 32'hf06f79a5;
        1573:    rdata = 32'h37b7b1bf;
        1574:    rdata = 32'he7170100;
        1575:    rdata = 32'h0713000e;
        1576:    rdata = 32'h86937b67;
        1577:    rdata = 32'hc31c0047;
        1578:    rdata = 32'h8693c354;
        1579:    rdata = 32'h07b10087;
        1580:    rdata = 32'hc75cc714;
        1581:    rdata = 32'h25b78082;
        1582:    rdata = 32'he5170100;
        1583:    rdata = 32'h0513000e;
        1584:    rdata = 32'hb1657a65;
        1585:    rdata = 32'h000ee797;
        1586:    rdata = 32'h7c078793;
        1587:    rdata = 32'hc3986741;
        1588:    rdata = 32'hc3d86711;
        1589:    rdata = 32'h00008082;
        1590:    rdata = 32'h00000000;
        1591:    rdata = 32'h00000000;
        1592:    rdata = 32'h00000000;
        1593:    rdata = 32'h00000000;
        1594:    rdata = 32'h00011876;
        1595:    rdata = 32'h00011886;
        1596:    rdata = 32'h00011896;
        1597:    rdata = 32'h000118b6;
        1598:    rdata = 32'h000118c4;
        1599:    rdata = 32'hffffecde;
        1600:    rdata = 32'hffffece4;
        1601:    rdata = 32'hffffecea;
        1602:    rdata = 32'hffffecf0;
        1603:    rdata = 32'hffffecfe;
        1604:    rdata = 32'hffffed06;
        1605:    rdata = 32'hffffed0e;
        1606:    rdata = 32'hffffed16;
        1607:    rdata = 32'hffffed1e;
        1608:    rdata = 32'hffffed24;
        1609:    rdata = 32'hffffed2a;
        1610:    rdata = 32'h0002c000;
        1611:    rdata = 32'h0003c000;
        1612:    rdata = 32'hc00002c0;
        1613:    rdata = 32'h02c00003;
        1614:    rdata = 32'h0003c000;
        1615:    rdata = 32'hc00002c0;
        1616:    rdata = 32'h02c00003;
        1617:    rdata = 32'h0003c000;
        1618:    rdata = 32'hc00002c0;
        1619:    rdata = 32'h02c00003;
        1620:    rdata = 32'h0003c000;
        1621:    rdata = 32'hc00002c0;
        1622:    rdata = 32'h02c00003;
        1623:    rdata = 32'h0003c000;
        1624:    rdata = 32'hc00002c0;
        1625:    rdata = 32'h02c00003;
        1626:    rdata = 32'h0003c000;
        1627:    rdata = 32'hc00002c0;
        1628:    rdata = 32'h02c00003;
        1629:    rdata = 32'h0003c000;
        1630:    rdata = 32'hc00002c0;
        1631:    rdata = 32'h02c00003;
        1632:    rdata = 32'h0003c000;
        1633:    rdata = 32'hc00002c0;
        1634:    rdata = 32'h02c00003;
        1635:    rdata = 32'h00042000;
        1636:    rdata = 32'h0020c000;
        1637:    rdata = 32'h200000c0;
        1638:    rdata = 32'h00000000;
        1639:    rdata = 32'h0008c000;
        1640:    rdata = 32'h200000c0;
        1641:    rdata = 32'h00000000;
        1642:    rdata = 32'h72616568;
        1643:    rdata = 32'h61656274;
        1644:    rdata = 32'h00000a74;
        1645:    rdata = 32'h706c6568;
        1646:    rdata = 32'h20202020;
        1647:    rdata = 32'h20202020;
        1648:    rdata = 32'h20202020;
        1649:    rdata = 32'h20202020;
        1650:    rdata = 32'h20202020;
        1651:    rdata = 32'h20202020;
        1652:    rdata = 32'h20202020;
        1653:    rdata = 32'h202d2020;
        1654:    rdata = 32'h6e697270;
        1655:    rdata = 32'h68742074;
        1656:    rdata = 32'h6d207369;
        1657:    rdata = 32'h61737365;
        1658:    rdata = 32'h720a6567;
        1659:    rdata = 32'h74657365;
        1660:    rdata = 32'h20202020;
        1661:    rdata = 32'h20202020;
        1662:    rdata = 32'h20202020;
        1663:    rdata = 32'h20202020;
        1664:    rdata = 32'h20202020;
        1665:    rdata = 32'h20202020;
        1666:    rdata = 32'h20202020;
        1667:    rdata = 32'h72202d20;
        1668:    rdata = 32'h74657365;
        1669:    rdata = 32'h636f7320;
        1670:    rdata = 32'h6e69700a;
        1671:    rdata = 32'h20202067;
        1672:    rdata = 32'h20202020;
        1673:    rdata = 32'h20202020;
        1674:    rdata = 32'h20202020;
        1675:    rdata = 32'h20202020;
        1676:    rdata = 32'h20202020;
        1677:    rdata = 32'h20202020;
        1678:    rdata = 32'h2d202020;
        1679:    rdata = 32'h6e657320;
        1680:    rdata = 32'h70222064;
        1681:    rdata = 32'h22676e69;
        1682:    rdata = 32'h206f7420;
        1683:    rdata = 32'h20656874;
        1684:    rdata = 32'h74736f68;
        1685:    rdata = 32'h7465730a;
        1686:    rdata = 32'h6970675f;
        1687:    rdata = 32'h69645f6f;
        1688:    rdata = 32'h74636572;
        1689:    rdata = 32'h206e6f69;
        1690:    rdata = 32'h6e69703c;
        1691:    rdata = 32'h695b203e;
        1692:    rdata = 32'h756f7c6e;
        1693:    rdata = 32'h2d205d74;
        1694:    rdata = 32'h74657320;
        1695:    rdata = 32'h69706720;
        1696:    rdata = 32'h6970206f;
        1697:    rdata = 32'h6964206e;
        1698:    rdata = 32'h74636572;
        1699:    rdata = 32'h0a6e6f69;
        1700:    rdata = 32'h5f746567;
        1701:    rdata = 32'h6f697067;
        1702:    rdata = 32'h7269645f;
        1703:    rdata = 32'h69746365;
        1704:    rdata = 32'h3c206e6f;
        1705:    rdata = 32'h3e6e6970;
        1706:    rdata = 32'h20202020;
        1707:    rdata = 32'h20202020;
        1708:    rdata = 32'h202d2020;
        1709:    rdata = 32'h20746567;
        1710:    rdata = 32'h6f697067;
        1711:    rdata = 32'h6e697020;
        1712:    rdata = 32'h72696420;
        1713:    rdata = 32'h69746365;
        1714:    rdata = 32'h730a6e6f;
        1715:    rdata = 32'h675f7465;
        1716:    rdata = 32'h206f6970;
        1717:    rdata = 32'h6e69703c;
        1718:    rdata = 32'h763c203e;
        1719:    rdata = 32'h65756c61;
        1720:    rdata = 32'h2020203e;
        1721:    rdata = 32'h20202020;
        1722:    rdata = 32'h20202020;
        1723:    rdata = 32'h73202d20;
        1724:    rdata = 32'h67207465;
        1725:    rdata = 32'h206f6970;
        1726:    rdata = 32'h0a6e6970;
        1727:    rdata = 32'h5f746567;
        1728:    rdata = 32'h6f697067;
        1729:    rdata = 32'h69703c20;
        1730:    rdata = 32'h20203e6e;
        1731:    rdata = 32'h20202020;
        1732:    rdata = 32'h20202020;
        1733:    rdata = 32'h20202020;
        1734:    rdata = 32'h20202020;
        1735:    rdata = 32'h202d2020;
        1736:    rdata = 32'h20746567;
        1737:    rdata = 32'h6f697067;
        1738:    rdata = 32'h6e697020;
        1739:    rdata = 32'h7465730a;
        1740:    rdata = 32'h6165685f;
        1741:    rdata = 32'h65627472;
        1742:    rdata = 32'h3c207461;
        1743:    rdata = 32'h69726570;
        1744:    rdata = 32'h5b20646f;
        1745:    rdata = 32'h3e5d736d;
        1746:    rdata = 32'h20202020;
        1747:    rdata = 32'h2d202020;
        1748:    rdata = 32'h74657320;
        1749:    rdata = 32'h61656820;
        1750:    rdata = 32'h65627472;
        1751:    rdata = 32'h720a7461;
        1752:    rdata = 32'h5f646165;
        1753:    rdata = 32'h7274616d;
        1754:    rdata = 32'h20207869;
        1755:    rdata = 32'h20202020;
        1756:    rdata = 32'h20202020;
        1757:    rdata = 32'h20202020;
        1758:    rdata = 32'h20202020;
        1759:    rdata = 32'h20202020;
        1760:    rdata = 32'h72202d20;
        1761:    rdata = 32'h20646165;
        1762:    rdata = 32'h7274616d;
        1763:    rdata = 32'h630a7869;
        1764:    rdata = 32'h62696c61;
        1765:    rdata = 32'h65746172;
        1766:    rdata = 32'h74616d5f;
        1767:    rdata = 32'h20786972;
        1768:    rdata = 32'h20202020;
        1769:    rdata = 32'h20202020;
        1770:    rdata = 32'h20202020;
        1771:    rdata = 32'h20202020;
        1772:    rdata = 32'h63202d20;
        1773:    rdata = 32'h62696c61;
        1774:    rdata = 32'h65746172;
        1775:    rdata = 32'h78697020;
        1776:    rdata = 32'h20736c65;
        1777:    rdata = 32'h7366666f;
        1778:    rdata = 32'h0a737465;
        1779:    rdata = 32'h00000000;
        1780:    rdata = 32'h6f727265;
        1781:    rdata = 32'h6f203a72;
        1782:    rdata = 32'h61726570;
        1783:    rdata = 32'h6e6f6974;
        1784:    rdata = 32'h746f6e20;
        1785:    rdata = 32'h70757320;
        1786:    rdata = 32'h74726f70;
        1787:    rdata = 32'h000a6465;
        1788:    rdata = 32'h676e6970;
        1789:    rdata = 32'h0000000a;
        1790:    rdata = 32'h6f727265;
        1791:    rdata = 32'h6d203a72;
        1792:    rdata = 32'h69737369;
        1793:    rdata = 32'h6120676e;
        1794:    rdata = 32'h6d756772;
        1795:    rdata = 32'h28746e65;
        1796:    rdata = 32'h000a2973;
        1797:    rdata = 32'h6f727265;
        1798:    rdata = 32'h69203a72;
        1799:    rdata = 32'h6c61766e;
        1800:    rdata = 32'h61206469;
        1801:    rdata = 32'h6d756772;
        1802:    rdata = 32'h28746e65;
        1803:    rdata = 32'h74202973;
        1804:    rdata = 32'h28657079;
        1805:    rdata = 32'h000a2973;
        1806:    rdata = 32'h00006e69;
        1807:    rdata = 32'h0074756f;
        1808:    rdata = 32'h6f727265;
        1809:    rdata = 32'h69203a72;
        1810:    rdata = 32'h6c61766e;
        1811:    rdata = 32'h64206469;
        1812:    rdata = 32'h63657269;
        1813:    rdata = 32'h6e6f6974;
        1814:    rdata = 32'h0000000a;
        1815:    rdata = 32'h6f727265;
        1816:    rdata = 32'h6d203a72;
        1817:    rdata = 32'h69737369;
        1818:    rdata = 32'h6120676e;
        1819:    rdata = 32'h6d756772;
        1820:    rdata = 32'h0a746e65;
        1821:    rdata = 32'h00000000;
        1822:    rdata = 32'h6f727265;
        1823:    rdata = 32'h69203a72;
        1824:    rdata = 32'h6c61766e;
        1825:    rdata = 32'h61206469;
        1826:    rdata = 32'h6d756772;
        1827:    rdata = 32'h20746e65;
        1828:    rdata = 32'h65707974;
        1829:    rdata = 32'h0000000a;
        1830:    rdata = 32'h64616572;
        1831:    rdata = 32'h5f74756f;
        1832:    rdata = 32'h656d6974;
        1833:    rdata = 32'h00000000;
        1834:    rdata = 32'h7366666f;
        1835:    rdata = 32'h63207465;
        1836:    rdata = 32'h62696c61;
        1837:    rdata = 32'h69746172;
        1838:    rdata = 32'h64206e6f;
        1839:    rdata = 32'h0a656e6f;
        1840:    rdata = 32'h00000000;
        1841:    rdata = 32'h696c6163;
        1842:    rdata = 32'h74617262;
        1843:    rdata = 32'h5f6e6f69;
        1844:    rdata = 32'h656d6974;
        1845:    rdata = 32'h00000000;
        1846:    rdata = 32'h0000203e;
        1847:    rdata = 32'h6f727265;
        1848:    rdata = 32'h75203a72;
        1849:    rdata = 32'h6365726e;
        1850:    rdata = 32'h696e676f;
        1851:    rdata = 32'h2064657a;
        1852:    rdata = 32'h6d6d6f63;
        1853:    rdata = 32'h3a646e61;
        1854:    rdata = 32'h00002220;
        1855:    rdata = 32'h65202e22;
        1856:    rdata = 32'h75636578;
        1857:    rdata = 32'h22206574;
        1858:    rdata = 32'h706c6568;
        1859:    rdata = 32'h6f742022;
        1860:    rdata = 32'h74656720;
        1861:    rdata = 32'h70757320;
        1862:    rdata = 32'h74726f70;
        1863:    rdata = 32'h63206465;
        1864:    rdata = 32'h616d6d6f;
        1865:    rdata = 32'h2073646e;
        1866:    rdata = 32'h7473696c;
        1867:    rdata = 32'h0000000a;
        1868:    rdata = 32'h6f727265;
        1869:    rdata = 32'h63203a72;
        1870:    rdata = 32'h616d6d6f;
        1871:    rdata = 32'h6620646e;
        1872:    rdata = 32'h656c6961;
        1873:    rdata = 32'h00000a64;
        1874:    rdata = 32'h706c6568;
        1875:    rdata = 32'h00000000;
        1876:    rdata = 32'h65736572;
        1877:    rdata = 32'h00000074;
        1878:    rdata = 32'h676e6970;
        1879:    rdata = 32'h00000000;
        1880:    rdata = 32'h5f746573;
        1881:    rdata = 32'h6f697067;
        1882:    rdata = 32'h7269645f;
        1883:    rdata = 32'h69746365;
        1884:    rdata = 32'h00006e6f;
        1885:    rdata = 32'h5f746567;
        1886:    rdata = 32'h6f697067;
        1887:    rdata = 32'h7269645f;
        1888:    rdata = 32'h69746365;
        1889:    rdata = 32'h00006e6f;
        1890:    rdata = 32'h5f746573;
        1891:    rdata = 32'h6f697067;
        1892:    rdata = 32'h00000000;
        1893:    rdata = 32'h5f746567;
        1894:    rdata = 32'h6f697067;
        1895:    rdata = 32'h00000000;
        1896:    rdata = 32'h5f746573;
        1897:    rdata = 32'h72616568;
        1898:    rdata = 32'h61656274;
        1899:    rdata = 32'h00000074;
        1900:    rdata = 32'h64616572;
        1901:    rdata = 32'h74616d5f;
        1902:    rdata = 32'h00786972;
        1903:    rdata = 32'h696c6163;
        1904:    rdata = 32'h74617262;
        1905:    rdata = 32'h616d5f65;
        1906:    rdata = 32'h78697274;
        1907:    rdata = 32'h00000000;
        1908:    rdata = 32'h6d6d6f63;
        1909:    rdata = 32'h5f646e61;
        1910:    rdata = 32'h65746e69;
        1911:    rdata = 32'h65727072;
        1912:    rdata = 32'h20726574;
        1913:    rdata = 32'h72617473;
        1914:    rdata = 32'h0a646574;
        1915:    rdata = 32'h00000000;
        1916:    rdata = 32'h0000203a;
        1917:    rdata = 32'h00002820;
        1918:    rdata = 32'h00203a29;
        1919:    rdata = 32'h6f636e69;
        1920:    rdata = 32'h63657272;
        1921:    rdata = 32'h61762074;
        1922:    rdata = 32'h2e65756c;
        1923:    rdata = 32'h79727420;
        1924:    rdata = 32'h61676120;
        1925:    rdata = 32'h000a6e69;
        default: rdata = 32'h00000000;
    endcase
end
endmodule
