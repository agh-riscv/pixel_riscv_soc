/**
 * Copyright (C) 2020  AGH University of Science and Technology
 *
 * This program is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with this program.  If not, see <https://www.gnu.org/licenses/>.
 */

module boot_mem (
    output logic [31:0] rdata,
    input logic [31:0] addr
);

/**
 * Module internal logic
 */

always_comb begin
    case (addr[13:2])
           0:    rdata = 32'h08c0006f;
           1:    rdata = 32'h0880006f;
           2:    rdata = 32'h0840006f;
           3:    rdata = 32'h0800006f;
           4:    rdata = 32'h07c0006f;
           5:    rdata = 32'h0780006f;
           6:    rdata = 32'h0740006f;
           7:    rdata = 32'h0700006f;
           8:    rdata = 32'h06c0006f;
           9:    rdata = 32'h0680006f;
          10:    rdata = 32'h0640006f;
          11:    rdata = 32'h0600006f;
          12:    rdata = 32'h05c0006f;
          13:    rdata = 32'h0580006f;
          14:    rdata = 32'h0540006f;
          15:    rdata = 32'h0500006f;
          16:    rdata = 32'h04c0006f;
          17:    rdata = 32'h0480006f;
          18:    rdata = 32'h0440006f;
          19:    rdata = 32'h0400006f;
          20:    rdata = 32'h03c0006f;
          21:    rdata = 32'h0380006f;
          22:    rdata = 32'h0340006f;
          23:    rdata = 32'h0300006f;
          24:    rdata = 32'h02c0006f;
          25:    rdata = 32'h0280006f;
          26:    rdata = 32'h0240006f;
          27:    rdata = 32'h0200006f;
          28:    rdata = 32'h01c0006f;
          29:    rdata = 32'h0180006f;
          30:    rdata = 32'h0140006f;
          31:    rdata = 32'h0100006f;
          32:    rdata = 32'h0100006f;
          33:    rdata = 32'h0080006f;
          34:    rdata = 32'h0040006f;
          35:    rdata = 32'h0000006f;
          36:    rdata = 32'h00000093;
          37:    rdata = 32'h00000113;
          38:    rdata = 32'h00000193;
          39:    rdata = 32'h00000213;
          40:    rdata = 32'h00000293;
          41:    rdata = 32'h00000313;
          42:    rdata = 32'h00000393;
          43:    rdata = 32'h00000413;
          44:    rdata = 32'h00000493;
          45:    rdata = 32'h00000513;
          46:    rdata = 32'h00000593;
          47:    rdata = 32'h00000613;
          48:    rdata = 32'h00000693;
          49:    rdata = 32'h00000713;
          50:    rdata = 32'h00000793;
          51:    rdata = 32'h00000813;
          52:    rdata = 32'h00000893;
          53:    rdata = 32'h00000913;
          54:    rdata = 32'h00000993;
          55:    rdata = 32'h00000a13;
          56:    rdata = 32'h00000a93;
          57:    rdata = 32'h00000b13;
          58:    rdata = 32'h00000b93;
          59:    rdata = 32'h00000c13;
          60:    rdata = 32'h00000c93;
          61:    rdata = 32'h00000d13;
          62:    rdata = 32'h00000d93;
          63:    rdata = 32'h00000e13;
          64:    rdata = 32'h00000e93;
          65:    rdata = 32'h00000f13;
          66:    rdata = 32'h00000f93;
          67:    rdata = 32'h00104117;
          68:    rdata = 32'hef410113;
          69:    rdata = 32'h00100297;
          70:    rdata = 32'heec28293;
          71:    rdata = 32'h00100317;
          72:    rdata = 32'hf3c30313;
          73:    rdata = 32'h0062d863;
          74:    rdata = 32'h0002a023;
          75:    rdata = 32'h00428293;
          76:    rdata = 32'hfe535ce3;
          77:    rdata = 32'h00001297;
          78:    rdata = 32'h8f428293;
          79:    rdata = 32'h00100317;
          80:    rdata = 32'hec430313;
          81:    rdata = 32'h00100397;
          82:    rdata = 32'hebc38393;
          83:    rdata = 32'h00735c63;
          84:    rdata = 32'h0002ae03;
          85:    rdata = 32'h01c32023;
          86:    rdata = 32'h00428293;
          87:    rdata = 32'h00430313;
          88:    rdata = 32'hfe7348e3;
          89:    rdata = 32'h00001297;
          90:    rdata = 32'h81028293;
          91:    rdata = 32'h00001317;
          92:    rdata = 32'h81830313;
          93:    rdata = 32'h0062da63;
          94:    rdata = 32'h0002a783;
          95:    rdata = 32'h000780e7;
          96:    rdata = 32'h00428293;
          97:    rdata = 32'hfe62cae3;
          98:    rdata = 32'h00000513;
          99:    rdata = 32'h00000593;
         100:    rdata = 32'h6e4000ef;
         101:    rdata = 32'h45857179;
         102:    rdata = 32'h00100517;
         103:    rdata = 32'he8c50513;
         104:    rdata = 32'hd422d606;
         105:    rdata = 32'hce4ed04a;
         106:    rdata = 32'hd226cc52;
         107:    rdata = 32'h458d2bbd;
         108:    rdata = 32'h00100517;
         109:    rdata = 32'he7450513;
         110:    rdata = 32'h44012b51;
         111:    rdata = 32'h00100917;
         112:    rdata = 32'he9490913;
         113:    rdata = 32'h00100997;
         114:    rdata = 32'he6098993;
         115:    rdata = 32'h854a4a11;
         116:    rdata = 32'h736329a1;
         117:    rdata = 32'h448102a4;
         118:    rdata = 32'h2bad854e;
         119:    rdata = 32'h97a6007c;
         120:    rdata = 32'h00a78023;
         121:    rdata = 32'h99e30485;
         122:    rdata = 32'h44b2ff44;
         123:    rdata = 32'h854a85a2;
         124:    rdata = 32'hc1042905;
         125:    rdata = 32'hbfe10411;
         126:    rdata = 32'h542250b2;
         127:    rdata = 32'h59025492;
         128:    rdata = 32'h4a6249f2;
         129:    rdata = 32'h80826145;
         130:    rdata = 32'hd4227179;
         131:    rdata = 32'hce4ed04a;
         132:    rdata = 32'hd606cc52;
         133:    rdata = 32'h4401d226;
         134:    rdata = 32'h00100917;
         135:    rdata = 32'he3890913;
         136:    rdata = 32'h00100997;
         137:    rdata = 32'he1898993;
         138:    rdata = 32'h854a4a11;
         139:    rdata = 32'h73632ef5;
         140:    rdata = 32'h448102a4;
         141:    rdata = 32'h2371854e;
         142:    rdata = 32'h97a6007c;
         143:    rdata = 32'h00a78023;
         144:    rdata = 32'h99e30485;
         145:    rdata = 32'h44b2ff44;
         146:    rdata = 32'h854a85a2;
         147:    rdata = 32'hc1042ed1;
         148:    rdata = 32'hbfe10411;
         149:    rdata = 32'h542250b2;
         150:    rdata = 32'h59025492;
         151:    rdata = 32'h4a6249f2;
         152:    rdata = 32'h80826145;
         153:    rdata = 32'hb73de111;
         154:    rdata = 32'h1141b745;
         155:    rdata = 32'h0613c422;
         156:    rdata = 32'h842a0640;
         157:    rdata = 32'h00100517;
         158:    rdata = 32'hdc450513;
         159:    rdata = 32'h2ba1c606;
         160:    rdata = 32'h852240b2;
         161:    rdata = 32'h01414422;
         162:    rdata = 32'h11418082;
         163:    rdata = 32'h842ac422;
         164:    rdata = 32'h00100517;
         165:    rdata = 32'hda850513;
         166:    rdata = 32'h237dc606;
         167:    rdata = 32'h852240b2;
         168:    rdata = 32'h01414422;
         169:    rdata = 32'h11418082;
         170:    rdata = 32'h842ac422;
         171:    rdata = 32'h00100517;
         172:    rdata = 32'hd8c50513;
         173:    rdata = 32'h2b49c606;
         174:    rdata = 32'h852240b2;
         175:    rdata = 32'h01414422;
         176:    rdata = 32'h418c8082;
         177:    rdata = 32'hcc221101;
         178:    rdata = 32'h0048842a;
         179:    rdata = 32'h2c19ce06;
         180:    rdata = 32'h0517004c;
         181:    rdata = 32'h05130010;
         182:    rdata = 32'h23bdd665;
         183:    rdata = 32'h852240f2;
         184:    rdata = 32'h61054462;
         185:    rdata = 32'h71758082;
         186:    rdata = 32'hc326c522;
         187:    rdata = 32'hdecec14a;
         188:    rdata = 32'hc706dcd2;
         189:    rdata = 32'h892e84aa;
         190:    rdata = 32'h00100417;
         191:    rdata = 32'hd4040413;
         192:    rdata = 32'h00000a17;
         193:    rdata = 32'h708a0a13;
         194:    rdata = 32'h00000997;
         195:    rdata = 32'h70498993;
         196:    rdata = 32'h852285ca;
         197:    rdata = 32'h85d22b15;
         198:    rdata = 32'h233d8522;
         199:    rdata = 32'h8526006c;
         200:    rdata = 32'h006837a9;
         201:    rdata = 32'he5092409;
         202:    rdata = 32'h852285ce;
         203:    rdata = 32'hb7cd2b31;
         204:    rdata = 32'h242d0068;
         205:    rdata = 32'h442a40ba;
         206:    rdata = 32'h490a449a;
         207:    rdata = 32'h5a6659f6;
         208:    rdata = 32'h80826149;
         209:    rdata = 32'h03000713;
         210:    rdata = 32'h00054783;
         211:    rdata = 32'h00e79463;
         212:    rdata = 32'hbfdd0505;
         213:    rdata = 32'h157de391;
         214:    rdata = 32'h47038082;
         215:    rdata = 32'h07930005;
         216:    rdata = 32'h136302d0;
         217:    rdata = 32'h050500f7;
         218:    rdata = 32'h47834725;
         219:    rdata = 32'h87930005;
         220:    rdata = 32'hf793fd07;
         221:    rdata = 32'h68630ff7;
         222:    rdata = 32'h478300f7;
         223:    rdata = 32'h05050015;
         224:    rdata = 32'h4505f7ed;
         225:    rdata = 32'h45018082;
         226:    rdata = 32'h05098082;
         227:    rdata = 32'h461546a5;
         228:    rdata = 32'h00054783;
         229:    rdata = 32'hfd078713;
         230:    rdata = 32'h0ff77713;
         231:    rdata = 32'h00e6fa63;
         232:    rdata = 32'hfdf7f793;
         233:    rdata = 32'hfbf78793;
         234:    rdata = 32'h0ff7f793;
         235:    rdata = 32'h00f66863;
         236:    rdata = 32'h00154783;
         237:    rdata = 32'hffe90505;
         238:    rdata = 32'h80824505;
         239:    rdata = 32'h80824501;
         240:    rdata = 32'hc70387aa;
         241:    rdata = 32'h05850005;
         242:    rdata = 32'h8fa30785;
         243:    rdata = 32'hfb75fee7;
         244:    rdata = 32'h87aa8082;
         245:    rdata = 32'h0007c683;
         246:    rdata = 32'h0785873e;
         247:    rdata = 32'hc783fee5;
         248:    rdata = 32'h05850005;
         249:    rdata = 32'h0fa30705;
         250:    rdata = 32'hfbf5fef7;
         251:    rdata = 32'h47838082;
         252:    rdata = 32'hc7030005;
         253:    rdata = 32'h87630005;
         254:    rdata = 32'h557d00e7;
         255:    rdata = 32'h00e7e963;
         256:    rdata = 32'h80824505;
         257:    rdata = 32'h0505c781;
         258:    rdata = 32'hb7d50585;
         259:    rdata = 32'h80824501;
         260:    rdata = 32'h450187aa;
         261:    rdata = 32'h00a78733;
         262:    rdata = 32'h00074703;
         263:    rdata = 32'h0505c319;
         264:    rdata = 32'h8082bfd5;
         265:    rdata = 32'h0c634789;
         266:    rdata = 32'h479102f6;
         267:    rdata = 32'h02f60d63;
         268:    rdata = 32'h47814705;
         269:    rdata = 32'h00e61463;
         270:    rdata = 32'h06400793;
         271:    rdata = 32'hcb8d4629;
         272:    rdata = 32'h02f5d733;
         273:    rdata = 32'h76930505;
         274:    rdata = 32'h86b30ff7;
         275:    rdata = 32'h071302f6;
         276:    rdata = 32'h0fa30307;
         277:    rdata = 32'hd7b3fee5;
         278:    rdata = 32'h8d9502c7;
         279:    rdata = 32'h6789b7cd;
         280:    rdata = 32'h71078793;
         281:    rdata = 32'hd7b7bfe1;
         282:    rdata = 32'h87933b9a;
         283:    rdata = 32'hb7f9a007;
         284:    rdata = 32'h00050023;
         285:    rdata = 32'h46058082;
         286:    rdata = 32'h1101b775;
         287:    rdata = 32'h4611cc22;
         288:    rdata = 32'h0048842a;
         289:    rdata = 32'h3f79ce06;
         290:    rdata = 32'h3d6d0048;
         291:    rdata = 32'h852285aa;
         292:    rdata = 32'h40f23f05;
         293:    rdata = 32'h61054462;
         294:    rdata = 32'h07938082;
         295:    rdata = 32'h06060300;
         296:    rdata = 32'h0ff67613;
         297:    rdata = 32'h00f50023;
         298:    rdata = 32'h07800793;
         299:    rdata = 32'h00f500a3;
         300:    rdata = 32'h87b24825;
         301:    rdata = 32'hf713c385;
         302:    rdata = 32'h069300f5;
         303:    rdata = 32'h64630577;
         304:    rdata = 32'h069300e8;
         305:    rdata = 32'h07330307;
         306:    rdata = 32'h00a300f5;
         307:    rdata = 32'h819100d7;
         308:    rdata = 32'hb7cd17fd;
         309:    rdata = 32'h01239532;
         310:    rdata = 32'h80820005;
         311:    rdata = 32'hbf754605;
         312:    rdata = 32'hbf654611;
         313:    rdata = 32'hcc221101;
         314:    rdata = 32'h842ace06;
         315:    rdata = 32'h0205d563;
         316:    rdata = 32'h02d00713;
         317:    rdata = 32'h00e50023;
         318:    rdata = 32'h40b005b3;
         319:    rdata = 32'h00484611;
         320:    rdata = 32'h00483715;
         321:    rdata = 32'h85aa3581;
         322:    rdata = 32'h00140513;
         323:    rdata = 32'h40f23d55;
         324:    rdata = 32'h61054462;
         325:    rdata = 32'h46118082;
         326:    rdata = 32'h37290048;
         327:    rdata = 32'h351d0048;
         328:    rdata = 32'h852285aa;
         329:    rdata = 32'h1141b7e5;
         330:    rdata = 32'hc606c422;
         331:    rdata = 32'h3535842a;
         332:    rdata = 32'h4703e115;
         333:    rdata = 32'h07930004;
         334:    rdata = 32'h1d630300;
         335:    rdata = 32'h470300f7;
         336:    rdata = 32'h07930014;
         337:    rdata = 32'h17630780;
         338:    rdata = 32'h852200f7;
         339:    rdata = 32'h40b24422;
         340:    rdata = 32'hbd250141;
         341:    rdata = 32'h442240b2;
         342:    rdata = 32'h80820141;
         343:    rdata = 32'hc4221141;
         344:    rdata = 32'h842ac606;
         345:    rdata = 32'h47833bdd;
         346:    rdata = 32'hc91d0004;
         347:    rdata = 32'h02d00693;
         348:    rdata = 32'h94634701;
         349:    rdata = 32'h872a00d7;
         350:    rdata = 32'h45010405;
         351:    rdata = 32'h46834629;
         352:    rdata = 32'hca810004;
         353:    rdata = 32'h02c507b3;
         354:    rdata = 32'hfd068513;
         355:    rdata = 32'h953e0405;
         356:    rdata = 32'hc319b7fd;
         357:    rdata = 32'h40a00533;
         358:    rdata = 32'h442240b2;
         359:    rdata = 32'h80820141;
         360:    rdata = 32'h03000713;
         361:    rdata = 32'h04e79663;
         362:    rdata = 32'h00144703;
         363:    rdata = 32'h07800793;
         364:    rdata = 32'h04f71063;
         365:    rdata = 32'h3bd18522;
         366:    rdata = 32'h0409cd05;
         367:    rdata = 32'h07134501;
         368:    rdata = 32'h06930600;
         369:    rdata = 32'h47830400;
         370:    rdata = 32'hd7f90004;
         371:    rdata = 32'h00f77a63;
         372:    rdata = 32'hfa978793;
         373:    rdata = 32'h0ff7f793;
         374:    rdata = 32'h8d5d0512;
         375:    rdata = 32'hb7e50405;
         376:    rdata = 32'h00f6f563;
         377:    rdata = 32'hfc978793;
         378:    rdata = 32'h8793b7f5;
         379:    rdata = 32'hb7ddfd07;
         380:    rdata = 32'hdeadc537;
         381:    rdata = 32'heef50513;
         382:    rdata = 32'h7793b745;
         383:    rdata = 32'h8793fdf5;
         384:    rdata = 32'hf793fbf7;
         385:    rdata = 32'h47650ff7;
         386:    rdata = 32'h00f77763;
         387:    rdata = 32'hfd050513;
         388:    rdata = 32'h00a53513;
         389:    rdata = 32'h45058082;
         390:    rdata = 32'hc10c8082;
         391:    rdata = 32'h8082c150;
         392:    rdata = 32'h99f14108;
         393:    rdata = 32'h8082952e;
         394:    rdata = 32'h80824148;
         395:    rdata = 32'h00458793;
         396:    rdata = 32'h8793c15c;
         397:    rdata = 32'hc51c0085;
         398:    rdata = 32'h00c58793;
         399:    rdata = 32'h8793c55c;
         400:    rdata = 32'hc91c0105;
         401:    rdata = 32'h01458793;
         402:    rdata = 32'h8793c95c;
         403:    rdata = 32'hc10c0185;
         404:    rdata = 32'h8793cd1c;
         405:    rdata = 32'h859301c5;
         406:    rdata = 32'hcd5c0205;
         407:    rdata = 32'h8082d10c;
         408:    rdata = 32'h8a05511c;
         409:    rdata = 32'h00b61633;
         410:    rdata = 32'h97b3439c;
         411:    rdata = 32'h8e5d48b7;
         412:    rdata = 32'hc390511c;
         413:    rdata = 32'h511c8082;
         414:    rdata = 32'h47854388;
         415:    rdata = 32'h00b797b3;
         416:    rdata = 32'h35338d7d;
         417:    rdata = 32'h808200a0;
         418:    rdata = 32'h4388455c;
         419:    rdata = 32'h97b34785;
         420:    rdata = 32'h8d7d00b7;
         421:    rdata = 32'h00a03533;
         422:    rdata = 32'h451c8082;
         423:    rdata = 32'h8e3d439c;
         424:    rdata = 32'h8e3d8e6d;
         425:    rdata = 32'hc390451c;
         426:    rdata = 32'h47858082;
         427:    rdata = 32'h00b61633;
         428:    rdata = 32'h00b795b3;
         429:    rdata = 32'h1141b7dd;
         430:    rdata = 32'hc226c422;
         431:    rdata = 32'h842ac606;
         432:    rdata = 32'h37d984ae;
         433:    rdata = 32'h00154613;
         434:    rdata = 32'h44228522;
         435:    rdata = 32'h85a640b2;
         436:    rdata = 32'h76134492;
         437:    rdata = 32'h01410ff6;
         438:    rdata = 32'h455cbfc9;
         439:    rdata = 32'h55134388;
         440:    rdata = 32'h80824915;
         441:    rdata = 32'h4388455c;
         442:    rdata = 32'h49055513;
         443:    rdata = 32'h11418082;
         444:    rdata = 32'h4601c226;
         445:    rdata = 32'h45bd84ae;
         446:    rdata = 32'hc606c422;
         447:    rdata = 32'h378d842a;
         448:    rdata = 32'h44228522;
         449:    rdata = 32'h862640b2;
         450:    rdata = 32'h45bd4492;
         451:    rdata = 32'hbf710141;
         452:    rdata = 32'h00458793;
         453:    rdata = 32'h8793c15c;
         454:    rdata = 32'hc10c0085;
         455:    rdata = 32'h8793c51c;
         456:    rdata = 32'h05c100c5;
         457:    rdata = 32'hc90cc55c;
         458:    rdata = 32'h41188082;
         459:    rdata = 32'h0015f793;
         460:    rdata = 32'h99f9430c;
         461:    rdata = 32'hc30c8ddd;
         462:    rdata = 32'h41188082;
         463:    rdata = 32'h97938985;
         464:    rdata = 32'h430c0015;
         465:    rdata = 32'h8ddd99f5;
         466:    rdata = 32'h8082c30c;
         467:    rdata = 32'h8023491c;
         468:    rdata = 32'h808200b7;
         469:    rdata = 32'h8023451c;
         470:    rdata = 32'h415c0007;
         471:    rdata = 32'h8b85439c;
         472:    rdata = 32'h455cdfed;
         473:    rdata = 32'h0007c503;
         474:    rdata = 32'h0ff57513;
         475:    rdata = 32'h451c8082;
         476:    rdata = 32'h00b78023;
         477:    rdata = 32'h439c415c;
         478:    rdata = 32'h4817d793;
         479:    rdata = 32'h455cffe5;
         480:    rdata = 32'h0007c783;
         481:    rdata = 32'h415c8082;
         482:    rdata = 32'h89054388;
         483:    rdata = 32'h415c8082;
         484:    rdata = 32'h55134388;
         485:    rdata = 32'h80824815;
         486:    rdata = 32'h00458793;
         487:    rdata = 32'h8793c15c;
         488:    rdata = 32'hc51c0085;
         489:    rdata = 32'h00c58793;
         490:    rdata = 32'h8793c55c;
         491:    rdata = 32'hc91c0105;
         492:    rdata = 32'hc10c47b1;
         493:    rdata = 32'h00f58823;
         494:    rdata = 32'he793419c;
         495:    rdata = 32'hc19c0017;
         496:    rdata = 32'h415c8082;
         497:    rdata = 32'h8b85439c;
         498:    rdata = 32'h455cdfed;
         499:    rdata = 32'h0007c503;
         500:    rdata = 32'h0ff57513;
         501:    rdata = 32'h11018082;
         502:    rdata = 32'hca26cc22;
         503:    rdata = 32'hc64ec84a;
         504:    rdata = 32'hc05ac256;
         505:    rdata = 32'hc452ce06;
         506:    rdata = 32'h892e84aa;
         507:    rdata = 32'h440189b2;
         508:    rdata = 32'h4b214aa9;
         509:    rdata = 32'h03345f63;
         510:    rdata = 32'h0a338526;
         511:    rdata = 32'h37d10089;
         512:    rdata = 32'h00aa0023;
         513:    rdata = 32'h01551f63;
         514:    rdata = 32'h000a0023;
         515:    rdata = 32'h40f24501;
         516:    rdata = 32'h44d24462;
         517:    rdata = 32'h49b24942;
         518:    rdata = 32'h4a924a22;
         519:    rdata = 32'h61054b02;
         520:    rdata = 32'h14638082;
         521:    rdata = 32'hc4010165;
         522:    rdata = 32'h04051479;
         523:    rdata = 32'h547db7e1;
         524:    rdata = 32'h4505bfed;
         525:    rdata = 32'h451cbfe9;
         526:    rdata = 32'h00b78023;
         527:    rdata = 32'h439c415c;
         528:    rdata = 32'h4817d793;
         529:    rdata = 32'h8082ffe5;
         530:    rdata = 32'hc4221141;
         531:    rdata = 32'hc606c226;
         532:    rdata = 32'h842e84aa;
         533:    rdata = 32'h00044583;
         534:    rdata = 32'h8526c589;
         535:    rdata = 32'h3fe10405;
         536:    rdata = 32'h40b2bfd5;
         537:    rdata = 32'h44924422;
         538:    rdata = 32'h80820141;
         539:    rdata = 32'h4388415c;
         540:    rdata = 32'h80828905;
         541:    rdata = 32'h05971141;
         542:    rdata = 32'h85930000;
         543:    rdata = 32'hf51710e5;
         544:    rdata = 32'h0513000f;
         545:    rdata = 32'hc6067ce5;
         546:    rdata = 32'h3c31c422;
         547:    rdata = 32'h000ff517;
         548:    rdata = 32'h77450513;
         549:    rdata = 32'h05973599;
         550:    rdata = 32'h85930000;
         551:    rdata = 32'he91d1025;
         552:    rdata = 32'h000ff517;
         553:    rdata = 32'h76050513;
         554:    rdata = 32'h842a3d35;
         555:    rdata = 32'h00000597;
         556:    rdata = 32'h10058593;
         557:    rdata = 32'h0597e509;
         558:    rdata = 32'h85930000;
         559:    rdata = 32'hf51710e5;
         560:    rdata = 32'h0513000f;
         561:    rdata = 32'h32c578e5;
         562:    rdata = 32'h3a698522;
         563:    rdata = 32'h00000597;
         564:    rdata = 32'h11058593;
         565:    rdata = 32'h000ff517;
         566:    rdata = 32'h77850513;
         567:    rdata = 32'h62c132e9;
         568:    rdata = 32'h305292f3;
         569:    rdata = 32'h00000597;
         570:    rdata = 32'h10c58593;
         571:    rdata = 32'h000ff517;
         572:    rdata = 32'h76050513;
         573:    rdata = 32'h45853a4d;
         574:    rdata = 32'h000ff517;
         575:    rdata = 32'h70850513;
         576:    rdata = 32'hf06f33fd;
         577:    rdata = 32'h40b277e0;
         578:    rdata = 32'h45014422;
         579:    rdata = 32'h80820141;
         580:    rdata = 32'h000ff797;
         581:    rdata = 32'h74078793;
         582:    rdata = 32'hc3986741;
         583:    rdata = 32'hc3d86711;
         584:    rdata = 32'h05b78082;
         585:    rdata = 32'hf5170100;
         586:    rdata = 32'h0513000f;
         587:    rdata = 32'hb9fd6da5;
         588:    rdata = 32'h010017b7;
         589:    rdata = 32'h000ff717;
         590:    rdata = 32'h6f070713;
         591:    rdata = 32'h00478693;
         592:    rdata = 32'h8693c354;
         593:    rdata = 32'hc31c0087;
         594:    rdata = 32'h8693c714;
         595:    rdata = 32'h07c100c7;
         596:    rdata = 32'hcb1cc754;
         597:    rdata = 32'h25b78082;
         598:    rdata = 32'hf5170100;
         599:    rdata = 32'h0513000f;
         600:    rdata = 32'hbd1d6de5;
         601:    rdata = 32'h00000000;
         602:    rdata = 32'h00000000;
         603:    rdata = 32'h00000000;
         604:    rdata = 32'h00000000;
         605:    rdata = 32'h00000910;
         606:    rdata = 32'h00000922;
         607:    rdata = 32'h00000930;
         608:    rdata = 32'h00000956;
         609:    rdata = 32'h746f6f62;
         610:    rdata = 32'h64616f6c;
         611:    rdata = 32'h73207265;
         612:    rdata = 32'h74726174;
         613:    rdata = 32'h000a6465;
         614:    rdata = 32'h65646f63;
         615:    rdata = 32'h64616f6c;
         616:    rdata = 32'h696b7320;
         617:    rdata = 32'h64657070;
         618:    rdata = 32'h0000000a;
         619:    rdata = 32'h65646f63;
         620:    rdata = 32'h64616f6c;
         621:    rdata = 32'h756f7320;
         622:    rdata = 32'h3a656372;
         623:    rdata = 32'h72617520;
         624:    rdata = 32'h00000a74;
         625:    rdata = 32'h65646f63;
         626:    rdata = 32'h64616f6c;
         627:    rdata = 32'h756f7320;
         628:    rdata = 32'h3a656372;
         629:    rdata = 32'h69707320;
         630:    rdata = 32'h0000000a;
         631:    rdata = 32'h65646f63;
         632:    rdata = 32'h64616f6c;
         633:    rdata = 32'h6e696620;
         634:    rdata = 32'h65687369;
         635:    rdata = 32'h00000a64;
         636:    rdata = 32'h746f6f62;
         637:    rdata = 32'h64616f6c;
         638:    rdata = 32'h66207265;
         639:    rdata = 32'h73696e69;
         640:    rdata = 32'h0a646568;
         641:    rdata = 32'h00000000;
         642:    rdata = 32'h0000203a;
         643:    rdata = 32'h6f636e69;
         644:    rdata = 32'h63657272;
         645:    rdata = 32'h61762074;
         646:    rdata = 32'h2e65756c;
         647:    rdata = 32'h79727420;
         648:    rdata = 32'h61676120;
         649:    rdata = 32'h000a6e69;
        default: rdata = 32'h00000000;
    endcase
end
endmodule
