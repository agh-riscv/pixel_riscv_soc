/**
 * Copyright (C) 2020  AGH University of Science and Technology
 *
 * This program is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with this program.  If not, see <https://www.gnu.org/licenses/>.
 */

module spi_mem (
    output logic [31:0] rdata,
    input logic [31:0] addr
);

/**
 * Module internal logic
 */

always_comb begin
    case (addr[13:2])
           0:    rdata = 32'h11b0106f;
           1:    rdata = 32'h0880006f;
           2:    rdata = 32'h0840006f;
           3:    rdata = 32'h0800006f;
           4:    rdata = 32'h07c0006f;
           5:    rdata = 32'h0780006f;
           6:    rdata = 32'h0740006f;
           7:    rdata = 32'h0700006f;
           8:    rdata = 32'h06c0006f;
           9:    rdata = 32'h0680006f;
          10:    rdata = 32'h0640006f;
          11:    rdata = 32'h0600006f;
          12:    rdata = 32'h05c0006f;
          13:    rdata = 32'h0580006f;
          14:    rdata = 32'h0540006f;
          15:    rdata = 32'h0500006f;
          16:    rdata = 32'h1450106f;
          17:    rdata = 32'h1930106f;
          18:    rdata = 32'h1e10106f;
          19:    rdata = 32'h22f0106f;
          20:    rdata = 32'h03c0006f;
          21:    rdata = 32'h0380006f;
          22:    rdata = 32'h0340006f;
          23:    rdata = 32'h0300006f;
          24:    rdata = 32'h02c0006f;
          25:    rdata = 32'h0280006f;
          26:    rdata = 32'h0240006f;
          27:    rdata = 32'h0200006f;
          28:    rdata = 32'h01c0006f;
          29:    rdata = 32'h0180006f;
          30:    rdata = 32'h0140006f;
          31:    rdata = 32'h0100006f;
          32:    rdata = 32'h0100006f;
          33:    rdata = 32'h0080006f;
          34:    rdata = 32'h0040006f;
          35:    rdata = 32'h0000006f;
          36:    rdata = 32'h00000093;
          37:    rdata = 32'h00000113;
          38:    rdata = 32'h00000193;
          39:    rdata = 32'h00000213;
          40:    rdata = 32'h00000293;
          41:    rdata = 32'h00000313;
          42:    rdata = 32'h00000393;
          43:    rdata = 32'h00000413;
          44:    rdata = 32'h00000493;
          45:    rdata = 32'h00000513;
          46:    rdata = 32'h00000593;
          47:    rdata = 32'h00000613;
          48:    rdata = 32'h00000693;
          49:    rdata = 32'h00000713;
          50:    rdata = 32'h00000793;
          51:    rdata = 32'h00000813;
          52:    rdata = 32'h00000893;
          53:    rdata = 32'h00000913;
          54:    rdata = 32'h00000993;
          55:    rdata = 32'h00000a13;
          56:    rdata = 32'h00000a93;
          57:    rdata = 32'h00000b13;
          58:    rdata = 32'h00000b93;
          59:    rdata = 32'h00000c13;
          60:    rdata = 32'h00000c93;
          61:    rdata = 32'h00000d13;
          62:    rdata = 32'h00000d93;
          63:    rdata = 32'h00000e13;
          64:    rdata = 32'h00000e93;
          65:    rdata = 32'h00000f13;
          66:    rdata = 32'h00000f93;
          67:    rdata = 32'h000f4117;
          68:    rdata = 32'hef410113;
          69:    rdata = 32'h000f0297;
          70:    rdata = 32'heec28293;
          71:    rdata = 32'h000f0317;
          72:    rdata = 32'hf2430313;
          73:    rdata = 32'h0062d863;
          74:    rdata = 32'h0002a023;
          75:    rdata = 32'h00428293;
          76:    rdata = 32'hfe535ce3;
          77:    rdata = 32'h00003297;
          78:    rdata = 32'hef428293;
          79:    rdata = 32'h000f0317;
          80:    rdata = 32'hec430313;
          81:    rdata = 32'h000f0397;
          82:    rdata = 32'hebc38393;
          83:    rdata = 32'h00735c63;
          84:    rdata = 32'h0002ae03;
          85:    rdata = 32'h01c32023;
          86:    rdata = 32'h00428293;
          87:    rdata = 32'h00430313;
          88:    rdata = 32'hfe7348e3;
          89:    rdata = 32'h00002297;
          90:    rdata = 32'h34028293;
          91:    rdata = 32'h00002317;
          92:    rdata = 32'h34c30313;
          93:    rdata = 32'h0062da63;
          94:    rdata = 32'h0002a783;
          95:    rdata = 32'h000780e7;
          96:    rdata = 32'h00428293;
          97:    rdata = 32'hfe62cae3;
          98:    rdata = 32'h00000513;
          99:    rdata = 32'h00000593;
         100:    rdata = 32'h296020ef;
         101:    rdata = 32'h35971141;
         102:    rdata = 32'h85930000;
         103:    rdata = 32'h051785a5;
         104:    rdata = 32'h0513000f;
         105:    rdata = 32'hc606e8e5;
         106:    rdata = 32'h61c010ef;
         107:    rdata = 32'h000f0517;
         108:    rdata = 32'he8c50513;
         109:    rdata = 32'h519010ef;
         110:    rdata = 32'h051740b2;
         111:    rdata = 32'h0513000f;
         112:    rdata = 32'h0141e7e5;
         113:    rdata = 32'h5390106f;
         114:    rdata = 32'h00003597;
         115:    rdata = 32'h83458593;
         116:    rdata = 32'h000f0517;
         117:    rdata = 32'he5c50513;
         118:    rdata = 32'h5ec0106f;
         119:    rdata = 32'h00003597;
         120:    rdata = 32'hb1858593;
         121:    rdata = 32'h000f0517;
         122:    rdata = 32'he4850513;
         123:    rdata = 32'h5d80106f;
         124:    rdata = 32'h00003597;
         125:    rdata = 32'hb2458593;
         126:    rdata = 32'h000f0517;
         127:    rdata = 32'he3450513;
         128:    rdata = 32'h5c40106f;
         129:    rdata = 32'h114141d8;
         130:    rdata = 32'hc422c606;
         131:    rdata = 32'hc04ac226;
         132:    rdata = 32'hc4634785;
         133:    rdata = 32'h359702e7;
         134:    rdata = 32'h85930000;
         135:    rdata = 32'h0517b065;
         136:    rdata = 32'h0513000f;
         137:    rdata = 32'h10efe0e5;
         138:    rdata = 32'h440559e0;
         139:    rdata = 32'h852240b2;
         140:    rdata = 32'h44924422;
         141:    rdata = 32'h01414902;
         142:    rdata = 32'h45808082;
         143:    rdata = 32'h146384ae;
         144:    rdata = 32'h559c00f4;
         145:    rdata = 32'h3597c791;
         146:    rdata = 32'h85930000;
         147:    rdata = 32'hbfc1af25;
         148:    rdata = 32'h02c58913;
         149:    rdata = 32'h3597854a;
         150:    rdata = 32'h85930000;
         151:    rdata = 32'h10efb065;
         152:    rdata = 32'hc50d2fa0;
         153:    rdata = 32'h00003597;
         154:    rdata = 32'hafc58593;
         155:    rdata = 32'h10ef854a;
         156:    rdata = 32'hcd012ea0;
         157:    rdata = 32'h00003597;
         158:    rdata = 32'haf058593;
         159:    rdata = 32'h000f0517;
         160:    rdata = 32'hdb050513;
         161:    rdata = 32'h540010ef;
         162:    rdata = 32'h4401b755;
         163:    rdata = 32'h00c4c583;
         164:    rdata = 32'h05178622;
         165:    rdata = 32'h0513000f;
         166:    rdata = 32'h10efd9e5;
         167:    rdata = 32'h44010370;
         168:    rdata = 32'h41dcb771;
         169:    rdata = 32'hc6061141;
         170:    rdata = 32'h02f04063;
         171:    rdata = 32'h00003597;
         172:    rdata = 32'had458593;
         173:    rdata = 32'h000f0517;
         174:    rdata = 32'hd7850513;
         175:    rdata = 32'h508010ef;
         176:    rdata = 32'h40b24505;
         177:    rdata = 32'h80820141;
         178:    rdata = 32'h47854598;
         179:    rdata = 32'h00f70763;
         180:    rdata = 32'h00003597;
         181:    rdata = 32'hacc58593;
         182:    rdata = 32'hc583bff1;
         183:    rdata = 32'h051700c5;
         184:    rdata = 32'h0513000f;
         185:    rdata = 32'h10efd525;
         186:    rdata = 32'h35977f80;
         187:    rdata = 32'h85930000;
         188:    rdata = 32'hc509a765;
         189:    rdata = 32'h00003597;
         190:    rdata = 32'ha6858593;
         191:    rdata = 32'h000f0517;
         192:    rdata = 32'hd3050513;
         193:    rdata = 32'h4c0010ef;
         194:    rdata = 32'h00003597;
         195:    rdata = 32'hab058593;
         196:    rdata = 32'h4b4010ef;
         197:    rdata = 32'hb7754501;
         198:    rdata = 32'h114141dc;
         199:    rdata = 32'h4705c606;
         200:    rdata = 32'h02f74063;
         201:    rdata = 32'h00003597;
         202:    rdata = 32'h9f858593;
         203:    rdata = 32'h000f0517;
         204:    rdata = 32'hd0050513;
         205:    rdata = 32'h490010ef;
         206:    rdata = 32'h40b24505;
         207:    rdata = 32'h80820141;
         208:    rdata = 32'h9563459c;
         209:    rdata = 32'h559800e7;
         210:    rdata = 32'h00f70763;
         211:    rdata = 32'h00003597;
         212:    rdata = 32'h9ec58593;
         213:    rdata = 32'h55d0bfe1;
         214:    rdata = 32'h00c5c583;
         215:    rdata = 32'h000f0517;
         216:    rdata = 32'hcd450513;
         217:    rdata = 32'h00c03633;
         218:    rdata = 32'h790010ef;
         219:    rdata = 32'hb7f14501;
         220:    rdata = 32'h110141dc;
         221:    rdata = 32'h4063ce06;
         222:    rdata = 32'h359702f0;
         223:    rdata = 32'h85930000;
         224:    rdata = 32'h0517a065;
         225:    rdata = 32'h0513000f;
         226:    rdata = 32'h10efcaa5;
         227:    rdata = 32'h450543a0;
         228:    rdata = 32'h610540f2;
         229:    rdata = 32'h45988082;
         230:    rdata = 32'h07634785;
         231:    rdata = 32'h359700f7;
         232:    rdata = 32'h85930000;
         233:    rdata = 32'hbff19fe5;
         234:    rdata = 32'h00c5c583;
         235:    rdata = 32'h000f0517;
         236:    rdata = 32'hc8450513;
         237:    rdata = 32'h752010ef;
         238:    rdata = 32'h006cc62a;
         239:    rdata = 32'h000f0517;
         240:    rdata = 32'hc7050513;
         241:    rdata = 32'h41e010ef;
         242:    rdata = 32'h00003597;
         243:    rdata = 32'h9f058593;
         244:    rdata = 32'h3f4010ef;
         245:    rdata = 32'hbf6d4501;
         246:    rdata = 32'h114141dc;
         247:    rdata = 32'hc422c606;
         248:    rdata = 32'h02f04163;
         249:    rdata = 32'h00003597;
         250:    rdata = 32'h99c58593;
         251:    rdata = 32'h000f0517;
         252:    rdata = 32'hc4050513;
         253:    rdata = 32'h3d0010ef;
         254:    rdata = 32'h40b24505;
         255:    rdata = 32'h01414422;
         256:    rdata = 32'h45988082;
         257:    rdata = 32'h842e4785;
         258:    rdata = 32'h00f70763;
         259:    rdata = 32'h00003597;
         260:    rdata = 32'h99058593;
         261:    rdata = 32'h45dcbfe1;
         262:    rdata = 32'h04f05d63;
         263:    rdata = 32'h00000597;
         264:    rdata = 32'hd7858593;
         265:    rdata = 32'h000f0517;
         266:    rdata = 32'hbdc50513;
         267:    rdata = 32'h4a0010ef;
         268:    rdata = 32'h67b1444c;
         269:    rdata = 32'h35078793;
         270:    rdata = 32'h02f585b3;
         271:    rdata = 32'h000f0517;
         272:    rdata = 32'hbfc50513;
         273:    rdata = 32'h10ef15fd;
         274:    rdata = 32'h05172690;
         275:    rdata = 32'h0513000f;
         276:    rdata = 32'h10efbee5;
         277:    rdata = 32'h05172b70;
         278:    rdata = 32'h0513000f;
         279:    rdata = 32'h10efbe25;
         280:    rdata = 32'h05172570;
         281:    rdata = 32'h0513000f;
         282:    rdata = 32'h10efb9e5;
         283:    rdata = 32'h45014400;
         284:    rdata = 32'h0517b769;
         285:    rdata = 32'h0513000f;
         286:    rdata = 32'h10efbc65;
         287:    rdata = 32'h05172470;
         288:    rdata = 32'h0513000f;
         289:    rdata = 32'h10efb825;
         290:    rdata = 32'hb7d54520;
         291:    rdata = 32'h110141d8;
         292:    rdata = 32'hcc22ce06;
         293:    rdata = 32'h4789ca26;
         294:    rdata = 32'h02e7c363;
         295:    rdata = 32'h00003597;
         296:    rdata = 32'h88058593;
         297:    rdata = 32'h000f0517;
         298:    rdata = 32'hb8850513;
         299:    rdata = 32'h318010ef;
         300:    rdata = 32'h40f24405;
         301:    rdata = 32'h44628522;
         302:    rdata = 32'h610544d2;
         303:    rdata = 32'h459c8082;
         304:    rdata = 32'h97634705;
         305:    rdata = 32'h558000e7;
         306:    rdata = 32'h45a4e401;
         307:    rdata = 32'h00f48763;
         308:    rdata = 32'h00003597;
         309:    rdata = 32'h86858593;
         310:    rdata = 32'hc783b7f1;
         311:    rdata = 32'h071302c5;
         312:    rdata = 32'h846302d0;
         313:    rdata = 32'h666306e7;
         314:    rdata = 32'h071302f7;
         315:    rdata = 32'h826302a0;
         316:    rdata = 32'h071306e7;
         317:    rdata = 32'h886302b0;
         318:    rdata = 32'h359702e7;
         319:    rdata = 32'h85930000;
         320:    rdata = 32'h05178de5;
         321:    rdata = 32'h0513000f;
         322:    rdata = 32'h10efb2a5;
         323:    rdata = 32'h84262ba0;
         324:    rdata = 32'h0713b74d;
         325:    rdata = 32'h92e302f0;
         326:    rdata = 32'h45f8fee7;
         327:    rdata = 32'h45dcc321;
         328:    rdata = 32'h02e7c7b3;
         329:    rdata = 32'h45dca021;
         330:    rdata = 32'h97ba45f8;
         331:    rdata = 32'h0517006c;
         332:    rdata = 32'h0513000f;
         333:    rdata = 32'hc63eafe5;
         334:    rdata = 32'h2aa010ef;
         335:    rdata = 32'h00003597;
         336:    rdata = 32'h87c58593;
         337:    rdata = 32'h280010ef;
         338:    rdata = 32'h45dcb7ad;
         339:    rdata = 32'h8f9945f8;
         340:    rdata = 32'h45dcbff1;
         341:    rdata = 32'h87b345f8;
         342:    rdata = 32'hbfc902e7;
         343:    rdata = 32'h00003597;
         344:    rdata = 32'h86058593;
         345:    rdata = 32'h41dcb781;
         346:    rdata = 32'hc6061141;
         347:    rdata = 32'hc226c422;
         348:    rdata = 32'h00f04e63;
         349:    rdata = 32'h00003597;
         350:    rdata = 32'h80c58593;
         351:    rdata = 32'h000f0517;
         352:    rdata = 32'hab050513;
         353:    rdata = 32'h240010ef;
         354:    rdata = 32'ha0ad4485;
         355:    rdata = 32'hc4914584;
         356:    rdata = 32'h00003597;
         357:    rdata = 32'h80c58593;
         358:    rdata = 32'h8413b7d5;
         359:    rdata = 32'h852200c5;
         360:    rdata = 32'h00003597;
         361:    rdata = 32'h85858593;
         362:    rdata = 32'h7b1000ef;
         363:    rdata = 32'hc11d4581;
         364:    rdata = 32'h00003597;
         365:    rdata = 32'h85458593;
         366:    rdata = 32'h00ef8522;
         367:    rdata = 32'h458579f0;
         368:    rdata = 32'h3597c911;
         369:    rdata = 32'h85930000;
         370:    rdata = 32'h852284e5;
         371:    rdata = 32'h78d000ef;
         372:    rdata = 32'h4589e905;
         373:    rdata = 32'h000f0517;
         374:    rdata = 32'ha4c50513;
         375:    rdata = 32'h6be000ef;
         376:    rdata = 32'h00003597;
         377:    rdata = 32'h85858593;
         378:    rdata = 32'h000f0517;
         379:    rdata = 32'ha4450513;
         380:    rdata = 32'h1d4010ef;
         381:    rdata = 32'h442240b2;
         382:    rdata = 32'h44928526;
         383:    rdata = 32'h80820141;
         384:    rdata = 32'h00003597;
         385:    rdata = 32'h81858593;
         386:    rdata = 32'h0113bf95;
         387:    rdata = 32'h4581df01;
         388:    rdata = 32'h000f0517;
         389:    rdata = 32'ha0450513;
         390:    rdata = 32'h20112623;
         391:    rdata = 32'h20812423;
         392:    rdata = 32'h20912223;
         393:    rdata = 32'h65e010ef;
         394:    rdata = 32'h000f0517;
         395:    rdata = 32'h9d850513;
         396:    rdata = 32'h25a010ef;
         397:    rdata = 32'h4685842a;
         398:    rdata = 32'h05974601;
         399:    rdata = 32'h8593000f;
         400:    rdata = 32'h850a9e65;
         401:    rdata = 32'h65a000ef;
         402:    rdata = 32'h000f0517;
         403:    rdata = 32'h9b850513;
         404:    rdata = 32'h23a010ef;
         405:    rdata = 32'h408505b3;
         406:    rdata = 32'h00002517;
         407:    rdata = 32'h7fc50513;
         408:    rdata = 32'h840a2391;
         409:    rdata = 32'h55030084;
         410:    rdata = 32'h04091c04;
         411:    rdata = 32'h1ce329e1;
         412:    rdata = 32'h2083fe94;
         413:    rdata = 32'h240320c1;
         414:    rdata = 32'h24832081;
         415:    rdata = 32'h01132041;
         416:    rdata = 32'h80822101;
         417:    rdata = 32'h45811141;
         418:    rdata = 32'h000f0517;
         419:    rdata = 32'h98c50513;
         420:    rdata = 32'hc422c606;
         421:    rdata = 32'h5ee010ef;
         422:    rdata = 32'h000f0517;
         423:    rdata = 32'h96850513;
         424:    rdata = 32'h1ea010ef;
         425:    rdata = 32'h0517842a;
         426:    rdata = 32'h0513000f;
         427:    rdata = 32'h00ef97a5;
         428:    rdata = 32'h05175ee0;
         429:    rdata = 32'h0513000f;
         430:    rdata = 32'h10ef94e5;
         431:    rdata = 32'h04331d00;
         432:    rdata = 32'h25974085;
         433:    rdata = 32'h85930000;
         434:    rdata = 32'h05177a25;
         435:    rdata = 32'h0513000f;
         436:    rdata = 32'h10ef9625;
         437:    rdata = 32'h85a20f20;
         438:    rdata = 32'h40b24422;
         439:    rdata = 32'h00002517;
         440:    rdata = 32'h7a450513;
         441:    rdata = 32'ha97d0141;
         442:    rdata = 32'hbf010113;
         443:    rdata = 32'h05174581;
         444:    rdata = 32'h0513000f;
         445:    rdata = 32'h26239325;
         446:    rdata = 32'h24234011;
         447:    rdata = 32'h2b714081;
         448:    rdata = 32'h00002617;
         449:    rdata = 32'hdf060613;
         450:    rdata = 32'h05174581;
         451:    rdata = 32'h0513000f;
         452:    rdata = 32'h00ef9165;
         453:    rdata = 32'h26175b00;
         454:    rdata = 32'h06130000;
         455:    rdata = 32'h4585fda6;
         456:    rdata = 32'h000f0517;
         457:    rdata = 32'h90050513;
         458:    rdata = 32'h59a000ef;
         459:    rdata = 32'h46014681;
         460:    rdata = 32'h000f0597;
         461:    rdata = 32'h8f058593;
         462:    rdata = 32'h2395850a;
         463:    rdata = 32'h05974605;
         464:    rdata = 32'h8593000f;
         465:    rdata = 32'h04088e25;
         466:    rdata = 32'h2b914681;
         467:    rdata = 32'h00002617;
         468:    rdata = 32'hda460613;
         469:    rdata = 32'h850a040c;
         470:    rdata = 32'h491010ef;
         471:    rdata = 32'h2617c911;
         472:    rdata = 32'h06130000;
         473:    rdata = 32'h0593f926;
         474:    rdata = 32'h04084001;
         475:    rdata = 32'h47d010ef;
         476:    rdata = 32'h00002597;
         477:    rdata = 32'h73458593;
         478:    rdata = 32'h0517842a;
         479:    rdata = 32'h0513000f;
         480:    rdata = 32'h10ef8b25;
         481:    rdata = 32'h25970420;
         482:    rdata = 32'h85930000;
         483:    rdata = 32'he40970e5;
         484:    rdata = 32'h00002597;
         485:    rdata = 32'h70c58593;
         486:    rdata = 32'h02c010ef;
         487:    rdata = 32'h40812403;
         488:    rdata = 32'h40c12083;
         489:    rdata = 32'h00002597;
         490:    rdata = 32'h61458593;
         491:    rdata = 32'h41010113;
         492:    rdata = 32'h0140106f;
         493:    rdata = 32'h2423714d;
         494:    rdata = 32'h22231481;
         495:    rdata = 32'h20231491;
         496:    rdata = 32'h2e231521;
         497:    rdata = 32'h2c231331;
         498:    rdata = 32'h2a231341;
         499:    rdata = 32'h28231351;
         500:    rdata = 32'h26231361;
         501:    rdata = 32'h842a1411;
         502:    rdata = 32'h00002a97;
         503:    rdata = 32'h6d4a8a93;
         504:    rdata = 32'h000f0497;
         505:    rdata = 32'h84c48493;
         506:    rdata = 32'h29174a35;
         507:    rdata = 32'h09130000;
         508:    rdata = 32'h2997cce9;
         509:    rdata = 32'h89930000;
         510:    rdata = 32'h2b177129;
         511:    rdata = 32'h0b130000;
         512:    rdata = 32'h85d66b6b;
         513:    rdata = 32'h00ef8526;
         514:    rdata = 32'h004c7bf0;
         515:    rdata = 32'h00ef8526;
         516:    rdata = 32'h00507770;
         517:    rdata = 32'h10a885a2;
         518:    rdata = 32'h57a62c71;
         519:    rdata = 32'hfefa63e3;
         520:    rdata = 32'h97ca078a;
         521:    rdata = 32'h97ca439c;
         522:    rdata = 32'h85228782;
         523:    rdata = 32'hbfd13a71;
         524:    rdata = 32'h326d8522;
         525:    rdata = 32'h8522b7f9;
         526:    rdata = 32'hb7e13a65;
         527:    rdata = 32'h852210ac;
         528:    rdata = 32'hd16132d1;
         529:    rdata = 32'h852685ce;
         530:    rdata = 32'h10aca8a9;
         531:    rdata = 32'h3c918522;
         532:    rdata = 32'h10acbfcd;
         533:    rdata = 32'h34c98522;
         534:    rdata = 32'h10acb7ed;
         535:    rdata = 32'h3e098522;
         536:    rdata = 32'h10acb7cd;
         537:    rdata = 32'h3e8d8522;
         538:    rdata = 32'h10acbfe9;
         539:    rdata = 32'h39398522;
         540:    rdata = 32'h10acbf49;
         541:    rdata = 32'h39c58522;
         542:    rdata = 32'h8522b769;
         543:    rdata = 32'hb7513379;
         544:    rdata = 32'h35098522;
         545:    rdata = 32'h8522bfbd;
         546:    rdata = 32'hbfa53585;
         547:    rdata = 32'h852685da;
         548:    rdata = 32'h735000ef;
         549:    rdata = 32'h00ef004c;
         550:    rdata = 32'h25977110;
         551:    rdata = 32'h85930000;
         552:    rdata = 32'h00ef6365;
         553:    rdata = 32'hbfb17230;
         554:    rdata = 32'h0713852e;
         555:    rdata = 32'h47830200;
         556:    rdata = 32'hc7890005;
         557:    rdata = 32'h00e79563;
         558:    rdata = 32'hbfd50505;
         559:    rdata = 32'h80824501;
         560:    rdata = 32'h00064783;
         561:    rdata = 32'h0df7f713;
         562:    rdata = 32'h0585c711;
         563:    rdata = 32'h8fa30605;
         564:    rdata = 32'hb7fdfef5;
         565:    rdata = 32'h00058023;
         566:    rdata = 32'hc7838082;
         567:    rdata = 32'hf7930005;
         568:    rdata = 32'hc3990df7;
         569:    rdata = 32'hbfd50585;
         570:    rdata = 32'hfff58513;
         571:    rdata = 32'h11018082;
         572:    rdata = 32'hc84acc22;
         573:    rdata = 32'hc256c452;
         574:    rdata = 32'hca26ce06;
         575:    rdata = 32'h892ac64e;
         576:    rdata = 32'h4a958432;
         577:    rdata = 32'h00860a13;
         578:    rdata = 32'hc6634044;
         579:    rdata = 32'h854a029a;
         580:    rdata = 32'h89aa3f61;
         581:    rdata = 32'h9593c10d;
         582:    rdata = 32'h05910054;
         583:    rdata = 32'h95d2862a;
         584:    rdata = 32'h3f79854a;
         585:    rdata = 32'h854a85ce;
         586:    rdata = 32'h405c3f4d;
         587:    rdata = 32'h00150593;
         588:    rdata = 32'hc05c0785;
         589:    rdata = 32'h40f2bfd1;
         590:    rdata = 32'h44d24462;
         591:    rdata = 32'h49b24942;
         592:    rdata = 32'h4a924a22;
         593:    rdata = 32'h80826105;
         594:    rdata = 32'hc2261141;
         595:    rdata = 32'h00c58493;
         596:    rdata = 32'h8526c422;
         597:    rdata = 32'h2597842e;
         598:    rdata = 32'h85930000;
         599:    rdata = 32'hc6065c65;
         600:    rdata = 32'h3f9000ef;
         601:    rdata = 32'h2023e919;
         602:    rdata = 32'h405c0004;
         603:    rdata = 32'h449240b2;
         604:    rdata = 32'hc05c17fd;
         605:    rdata = 32'h01414422;
         606:    rdata = 32'h25978082;
         607:    rdata = 32'h85930000;
         608:    rdata = 32'h85265aa5;
         609:    rdata = 32'h3d5000ef;
         610:    rdata = 32'hc5694785;
         611:    rdata = 32'h00002597;
         612:    rdata = 32'h5a058593;
         613:    rdata = 32'h00ef8526;
         614:    rdata = 32'h47893c30;
         615:    rdata = 32'h2597cd45;
         616:    rdata = 32'h85930000;
         617:    rdata = 32'h85265965;
         618:    rdata = 32'h3b1000ef;
         619:    rdata = 32'hc15d478d;
         620:    rdata = 32'h00002597;
         621:    rdata = 32'h59858593;
         622:    rdata = 32'h00ef8526;
         623:    rdata = 32'h479139f0;
         624:    rdata = 32'h2597c951;
         625:    rdata = 32'h85930000;
         626:    rdata = 32'h852659a5;
         627:    rdata = 32'h38d000ef;
         628:    rdata = 32'hc1494795;
         629:    rdata = 32'h00002597;
         630:    rdata = 32'h59458593;
         631:    rdata = 32'h00ef8526;
         632:    rdata = 32'h479937b0;
         633:    rdata = 32'h2597c925;
         634:    rdata = 32'h85930000;
         635:    rdata = 32'h852658e5;
         636:    rdata = 32'h369000ef;
         637:    rdata = 32'hcd39479d;
         638:    rdata = 32'h00002597;
         639:    rdata = 32'h58c58593;
         640:    rdata = 32'h00ef8526;
         641:    rdata = 32'h47a13570;
         642:    rdata = 32'h2597c531;
         643:    rdata = 32'h85930000;
         644:    rdata = 32'h85265865;
         645:    rdata = 32'h345000ef;
         646:    rdata = 32'hcd0d47a5;
         647:    rdata = 32'h00002597;
         648:    rdata = 32'h58c58593;
         649:    rdata = 32'h00ef8526;
         650:    rdata = 32'h47a93330;
         651:    rdata = 32'h2597c505;
         652:    rdata = 32'h85930000;
         653:    rdata = 32'h85265865;
         654:    rdata = 32'h321000ef;
         655:    rdata = 32'hc91947ad;
         656:    rdata = 32'h00002597;
         657:    rdata = 32'h58858593;
         658:    rdata = 32'h00ef8526;
         659:    rdata = 32'h47b130f0;
         660:    rdata = 32'h47b5c111;
         661:    rdata = 32'hbf11c01c;
         662:    rdata = 32'hcc221101;
         663:    rdata = 32'hc64ec84a;
         664:    rdata = 32'hce06c452;
         665:    rdata = 32'h892eca26;
         666:    rdata = 32'h00c58413;
         667:    rdata = 32'h4a054981;
         668:    rdata = 32'h00492783;
         669:    rdata = 32'h02f9d863;
         670:    rdata = 32'h02040493;
         671:    rdata = 32'h09858526;
         672:    rdata = 32'h411000ef;
         673:    rdata = 32'h2e23c909;
         674:    rdata = 32'h8526ff44;
         675:    rdata = 32'h43b000ef;
         676:    rdata = 32'h8426c008;
         677:    rdata = 32'h2e23bff1;
         678:    rdata = 32'h85a6fe04;
         679:    rdata = 32'h00ef8522;
         680:    rdata = 32'hbfc528d0;
         681:    rdata = 32'h446240f2;
         682:    rdata = 32'h494244d2;
         683:    rdata = 32'h4a2249b2;
         684:    rdata = 32'h80826105;
         685:    rdata = 32'hc6061141;
         686:    rdata = 32'hc226c422;
         687:    rdata = 32'h842ac04a;
         688:    rdata = 32'h893284ae;
         689:    rdata = 32'h00052223;
         690:    rdata = 32'h0c000613;
         691:    rdata = 32'h05214581;
         692:    rdata = 32'h03d010ef;
         693:    rdata = 32'h85ca8622;
         694:    rdata = 32'h3d118526;
         695:    rdata = 32'heb91405c;
         696:    rdata = 32'hc01c47b9;
         697:    rdata = 32'h852240b2;
         698:    rdata = 32'h44924422;
         699:    rdata = 32'h01414902;
         700:    rdata = 32'h85a28082;
         701:    rdata = 32'h3d898526;
         702:    rdata = 32'h852685a2;
         703:    rdata = 32'hb7dd3fb1;
         704:    rdata = 32'h85aa7119;
         705:    rdata = 32'hde860068;
         706:    rdata = 32'h223000ef;
         707:    rdata = 32'h00002597;
         708:    rdata = 32'h2ac58593;
         709:    rdata = 32'h00ef0068;
         710:    rdata = 32'h006c2270;
         711:    rdata = 32'h000ef517;
         712:    rdata = 32'h51050513;
         713:    rdata = 32'h4a1000ef;
         714:    rdata = 32'h610950f6;
         715:    rdata = 32'h11018082;
         716:    rdata = 32'h004885aa;
         717:    rdata = 32'h00efce06;
         718:    rdata = 32'h00482af0;
         719:    rdata = 32'h40f237d1;
         720:    rdata = 32'h80826105;
         721:    rdata = 32'h85aa1101;
         722:    rdata = 32'hce060048;
         723:    rdata = 32'h2ff000ef;
         724:    rdata = 32'h377d0048;
         725:    rdata = 32'h610540f2;
         726:    rdata = 32'h71198082;
         727:    rdata = 32'h842edca2;
         728:    rdata = 32'h006885aa;
         729:    rdata = 32'h00efde86;
         730:    rdata = 32'h25971c50;
         731:    rdata = 32'h85930000;
         732:    rdata = 32'h00684965;
         733:    rdata = 32'h1c9000ef;
         734:    rdata = 32'h006885a2;
         735:    rdata = 32'h1c1000ef;
         736:    rdata = 32'h00002597;
         737:    rdata = 32'h23858593;
         738:    rdata = 32'h00ef0068;
         739:    rdata = 32'h006c1b30;
         740:    rdata = 32'h000ef517;
         741:    rdata = 32'h49c50513;
         742:    rdata = 32'h42d000ef;
         743:    rdata = 32'h546650f6;
         744:    rdata = 32'h80826109;
         745:    rdata = 32'hcc221101;
         746:    rdata = 32'h0048842a;
         747:    rdata = 32'h00efce06;
         748:    rdata = 32'h004c2370;
         749:    rdata = 32'h37558522;
         750:    rdata = 32'h446240f2;
         751:    rdata = 32'h80826105;
         752:    rdata = 32'hcc221101;
         753:    rdata = 32'h0048842a;
         754:    rdata = 32'h00efce06;
         755:    rdata = 32'h004c2810;
         756:    rdata = 32'h37618522;
         757:    rdata = 32'h446240f2;
         758:    rdata = 32'h80826105;
         759:    rdata = 32'hdaa67119;
         760:    rdata = 32'h85aa84ae;
         761:    rdata = 32'hde860068;
         762:    rdata = 32'h8432dca2;
         763:    rdata = 32'h13f000ef;
         764:    rdata = 32'h00002597;
         765:    rdata = 32'h41458593;
         766:    rdata = 32'h00ef0068;
         767:    rdata = 32'h85a61430;
         768:    rdata = 32'h00ef0068;
         769:    rdata = 32'h259713b0;
         770:    rdata = 32'h85930000;
         771:    rdata = 32'h00684025;
         772:    rdata = 32'h12d000ef;
         773:    rdata = 32'h006885a2;
         774:    rdata = 32'h125000ef;
         775:    rdata = 32'h00002597;
         776:    rdata = 32'h19c58593;
         777:    rdata = 32'h00ef0068;
         778:    rdata = 32'h006c1170;
         779:    rdata = 32'h000ef517;
         780:    rdata = 32'h40050513;
         781:    rdata = 32'h391000ef;
         782:    rdata = 32'h546650f6;
         783:    rdata = 32'h610954d6;
         784:    rdata = 32'h71798082;
         785:    rdata = 32'h842ad422;
         786:    rdata = 32'hd6060028;
         787:    rdata = 32'h84b2d226;
         788:    rdata = 32'h1fb000ef;
         789:    rdata = 32'h084885a6;
         790:    rdata = 32'h18d000ef;
         791:    rdata = 32'h002c0850;
         792:    rdata = 32'h3fad8522;
         793:    rdata = 32'h542250b2;
         794:    rdata = 32'h61455492;
         795:    rdata = 32'h71798082;
         796:    rdata = 32'h842ad422;
         797:    rdata = 32'hd6060028;
         798:    rdata = 32'h84b2d226;
         799:    rdata = 32'h1cf000ef;
         800:    rdata = 32'h084885a6;
         801:    rdata = 32'h1c7000ef;
         802:    rdata = 32'h002c0850;
         803:    rdata = 32'h37b98522;
         804:    rdata = 32'h542250b2;
         805:    rdata = 32'h61455492;
         806:    rdata = 32'ha8898082;
         807:    rdata = 32'h1101abf5;
         808:    rdata = 32'hce06cc22;
         809:    rdata = 32'hc699842a;
         810:    rdata = 32'hc632852e;
         811:    rdata = 32'h285dc42e;
         812:    rdata = 32'h45a24632;
         813:    rdata = 32'h2ce98522;
         814:    rdata = 32'h852240f2;
         815:    rdata = 32'h61054462;
         816:    rdata = 32'habd18082;
         817:    rdata = 32'hc4221141;
         818:    rdata = 32'h842ac606;
         819:    rdata = 32'h85222181;
         820:    rdata = 32'h40b24422;
         821:    rdata = 32'ha8d90141;
         822:    rdata = 32'hc4221141;
         823:    rdata = 32'h842ac606;
         824:    rdata = 32'h85222b5d;
         825:    rdata = 32'h40b24422;
         826:    rdata = 32'ha0c90141;
         827:    rdata = 32'hc6061141;
         828:    rdata = 32'h4705c10c;
         829:    rdata = 32'h02e58563;
         830:    rdata = 32'h8b634709;
         831:    rdata = 32'he1a502e5;
         832:    rdata = 32'h000ef517;
         833:    rdata = 32'h31450513;
         834:    rdata = 32'h725000ef;
         835:    rdata = 32'h40b24581;
         836:    rdata = 32'h000ef517;
         837:    rdata = 32'h30450513;
         838:    rdata = 32'h006f0141;
         839:    rdata = 32'h458171f0;
         840:    rdata = 32'h000ef517;
         841:    rdata = 32'h2f450513;
         842:    rdata = 32'h705000ef;
         843:    rdata = 32'hb7c54585;
         844:    rdata = 32'hf5174585;
         845:    rdata = 32'h0513000e;
         846:    rdata = 32'h00ef2e25;
         847:    rdata = 32'h45856f30;
         848:    rdata = 32'h000ef517;
         849:    rdata = 32'h2d450513;
         850:    rdata = 32'h6f1000ef;
         851:    rdata = 32'h458140b2;
         852:    rdata = 32'h000ef517;
         853:    rdata = 32'h2c450513;
         854:    rdata = 32'h006f0141;
         855:    rdata = 32'h40b27030;
         856:    rdata = 32'h80820141;
         857:    rdata = 32'h11414118;
         858:    rdata = 32'h4785c606;
         859:    rdata = 32'h02e7e063;
         860:    rdata = 32'h000ef517;
         861:    rdata = 32'h2b850513;
         862:    rdata = 32'h720000ef;
         863:    rdata = 32'hf51740b2;
         864:    rdata = 32'h0513000e;
         865:    rdata = 32'h01412965;
         866:    rdata = 32'h0fe0106f;
         867:    rdata = 32'hf51745a1;
         868:    rdata = 32'h0513000e;
         869:    rdata = 32'h00ef2865;
         870:    rdata = 32'h40b26c70;
         871:    rdata = 32'hf5174581;
         872:    rdata = 32'h0513000e;
         873:    rdata = 32'h01412765;
         874:    rdata = 32'h6b50006f;
         875:    rdata = 32'h11414118;
         876:    rdata = 32'h4785c606;
         877:    rdata = 32'h02e7e063;
         878:    rdata = 32'h000ef517;
         879:    rdata = 32'h27050513;
         880:    rdata = 32'h6c2000ef;
         881:    rdata = 32'hf51740b2;
         882:    rdata = 32'h0513000e;
         883:    rdata = 32'h014124e5;
         884:    rdata = 32'h0b60106f;
         885:    rdata = 32'h02000593;
         886:    rdata = 32'h000ef517;
         887:    rdata = 32'h23c50513;
         888:    rdata = 32'h67d000ef;
         889:    rdata = 32'h458140b2;
         890:    rdata = 32'h000ef517;
         891:    rdata = 32'h22c50513;
         892:    rdata = 32'h006f0141;
         893:    rdata = 32'h419c66b0;
         894:    rdata = 32'hd4227179;
         895:    rdata = 32'hd226d606;
         896:    rdata = 32'hce4ed04a;
         897:    rdata = 32'hca56cc52;
         898:    rdata = 32'hc65ec85a;
         899:    rdata = 32'h842ac462;
         900:    rdata = 32'h4581eba5;
         901:    rdata = 32'h000ef517;
         902:    rdata = 32'h21450513;
         903:    rdata = 32'hf5172d29;
         904:    rdata = 32'h0513000e;
         905:    rdata = 32'h10ef1f65;
         906:    rdata = 32'hf4970600;
         907:    rdata = 32'h8493000e;
         908:    rdata = 32'h85261ea4;
         909:    rdata = 32'h05e010ef;
         910:    rdata = 32'h449ddd6d;
         911:    rdata = 32'h000ef917;
         912:    rdata = 32'h1d890913;
         913:    rdata = 32'h854a59fd;
         914:    rdata = 32'h03e010ef;
         915:    rdata = 32'h10ef854a;
         916:    rdata = 32'hdd6d0440;
         917:    rdata = 32'h00649593;
         918:    rdata = 32'h854a95a2;
         919:    rdata = 32'h00ef14fd;
         920:    rdata = 32'h92e363b0;
         921:    rdata = 32'h50b2ff34;
         922:    rdata = 32'h54228522;
         923:    rdata = 32'h59025492;
         924:    rdata = 32'h4a6249f2;
         925:    rdata = 32'h4b424ad2;
         926:    rdata = 32'h4c224bb2;
         927:    rdata = 32'h80826145;
         928:    rdata = 32'h9e634705;
         929:    rdata = 32'h458506e7;
         930:    rdata = 32'h000ef517;
         931:    rdata = 32'h1a050513;
         932:    rdata = 32'h449d235d;
         933:    rdata = 32'h000ef997;
         934:    rdata = 32'h18098993;
         935:    rdata = 32'h0b934b05;
         936:    rdata = 32'h5afd0200;
         937:    rdata = 32'h00649a13;
         938:    rdata = 32'h493d9a22;
         939:    rdata = 32'h00ef854e;
         940:    rdata = 32'h16335e50;
         941:    rdata = 32'h0642012b;
         942:    rdata = 32'h48138641;
         943:    rdata = 32'h8752fff6;
         944:    rdata = 32'h15b34681;
         945:    rdata = 32'h8de900db;
         946:    rdata = 32'h00071783;
         947:    rdata = 32'h8fd1c595;
         948:    rdata = 32'h00f71023;
         949:    rdata = 32'h07090685;
         950:    rdata = 32'hff7695e3;
         951:    rdata = 32'h00ef854e;
         952:    rdata = 32'hdd6d7b50;
         953:    rdata = 32'h197d854e;
         954:    rdata = 32'h79f000ef;
         955:    rdata = 32'hfd5910e3;
         956:    rdata = 32'h99e314fd;
         957:    rdata = 32'hbf85fb54;
         958:    rdata = 32'h00f877b3;
         959:    rdata = 32'h89b2bfd1;
         960:    rdata = 32'hc2114589;
         961:    rdata = 32'hf5174591;
         962:    rdata = 32'h0513000e;
         963:    rdata = 32'h00ef10e5;
         964:    rdata = 32'h491d54f0;
         965:    rdata = 32'h000ef497;
         966:    rdata = 32'h10048493;
         967:    rdata = 32'h0c134b85;
         968:    rdata = 32'h5b7d0200;
         969:    rdata = 32'h00691a93;
         970:    rdata = 32'h4a3d9aa2;
         971:    rdata = 32'h00ef8526;
         972:    rdata = 32'h96335650;
         973:    rdata = 32'h0642014b;
         974:    rdata = 32'h48138641;
         975:    rdata = 32'h8756fff6;
         976:    rdata = 32'h95b34681;
         977:    rdata = 32'h8de900db;
         978:    rdata = 32'h00071783;
         979:    rdata = 32'h8fd1c98d;
         980:    rdata = 32'h00f71023;
         981:    rdata = 32'h07090685;
         982:    rdata = 32'hff8695e3;
         983:    rdata = 32'h02099463;
         984:    rdata = 32'h8526458d;
         985:    rdata = 32'h4f9000ef;
         986:    rdata = 32'h85264589;
         987:    rdata = 32'h00ef1a7d;
         988:    rdata = 32'h1de34ef0;
         989:    rdata = 32'h197dfb6a;
         990:    rdata = 32'hfb6916e3;
         991:    rdata = 32'h77b3b5ed;
         992:    rdata = 32'hb7f900f8;
         993:    rdata = 32'h85264595;
         994:    rdata = 32'h4d5000ef;
         995:    rdata = 32'hbff14591;
         996:    rdata = 32'hc4221141;
         997:    rdata = 32'h842ac606;
         998:    rdata = 32'h40b23db9;
         999:    rdata = 32'h44228522;
        1000:    rdata = 32'h80820141;
        1001:    rdata = 32'h7159411c;
        1002:    rdata = 32'hd2a6d4a2;
        1003:    rdata = 32'hd0cad686;
        1004:    rdata = 32'hccd2cece;
        1005:    rdata = 32'hc8dacad6;
        1006:    rdata = 32'h842ec6de;
        1007:    rdata = 32'hefbd84b2;
        1008:    rdata = 32'h892a878a;
        1009:    rdata = 32'h902385be;
        1010:    rdata = 32'h00980097;
        1011:    rdata = 32'h9ce30789;
        1012:    rdata = 32'hf517fee7;
        1013:    rdata = 32'h0513000e;
        1014:    rdata = 32'h00ef0425;
        1015:    rdata = 32'h25834af0;
        1016:    rdata = 32'h86220009;
        1017:    rdata = 32'h000ef517;
        1018:    rdata = 32'h04450513;
        1019:    rdata = 32'hf51721a9;
        1020:    rdata = 32'h0513000e;
        1021:    rdata = 32'h00ef0265;
        1022:    rdata = 32'hf4176910;
        1023:    rdata = 32'h0413000e;
        1024:    rdata = 32'h852201a4;
        1025:    rdata = 32'h68f000ef;
        1026:    rdata = 32'h4421dd6d;
        1027:    rdata = 32'h000ef497;
        1028:    rdata = 32'h00848493;
        1029:    rdata = 32'h00ef8526;
        1030:    rdata = 32'h85266710;
        1031:    rdata = 32'h677000ef;
        1032:    rdata = 32'h147ddd6d;
        1033:    rdata = 32'h50b6f865;
        1034:    rdata = 32'h54965426;
        1035:    rdata = 32'h49f65906;
        1036:    rdata = 32'h4ad64a66;
        1037:    rdata = 32'h4bb64b46;
        1038:    rdata = 32'h80826165;
        1039:    rdata = 32'h4a214705;
        1040:    rdata = 32'h04e78a63;
        1041:    rdata = 32'h0b134a85;
        1042:    rdata = 32'hf9170200;
        1043:    rdata = 32'h0913000e;
        1044:    rdata = 32'h5bfdfca9;
        1045:    rdata = 32'hd6b349bd;
        1046:    rdata = 32'h8a854134;
        1047:    rdata = 32'h45814781;
        1048:    rdata = 32'h00fa9733;
        1049:    rdata = 32'h8dd9cad1;
        1050:    rdata = 32'h9be30785;
        1051:    rdata = 32'h854aff67;
        1052:    rdata = 32'h413000ef;
        1053:    rdata = 32'h458de451;
        1054:    rdata = 32'h00ef854a;
        1055:    rdata = 32'h45893e30;
        1056:    rdata = 32'h19fd854a;
        1057:    rdata = 32'h3d9000ef;
        1058:    rdata = 32'hfd7997e3;
        1059:    rdata = 32'h13e31a7d;
        1060:    rdata = 32'hbf51fc0a;
        1061:    rdata = 32'hf517862e;
        1062:    rdata = 32'h0513000e;
        1063:    rdata = 32'h4585f925;
        1064:    rdata = 32'h49212e59;
        1065:    rdata = 32'h0a934a05;
        1066:    rdata = 32'hf9970200;
        1067:    rdata = 32'h8993000e;
        1068:    rdata = 32'h5b7df6a9;
        1069:    rdata = 32'hd6b3443d;
        1070:    rdata = 32'h8a854084;
        1071:    rdata = 32'h45814781;
        1072:    rdata = 32'h00fa1733;
        1073:    rdata = 32'h8dd9c695;
        1074:    rdata = 32'h9be30785;
        1075:    rdata = 32'h854eff57;
        1076:    rdata = 32'h3b3000ef;
        1077:    rdata = 32'h00ef854e;
        1078:    rdata = 32'hdd6d5bd0;
        1079:    rdata = 32'h147d854e;
        1080:    rdata = 32'h5a7000ef;
        1081:    rdata = 32'hfd6419e3;
        1082:    rdata = 32'h15e3197d;
        1083:    rdata = 32'hbf25fc09;
        1084:    rdata = 32'hfff74713;
        1085:    rdata = 32'hbfc98df9;
        1086:    rdata = 32'hfff74713;
        1087:    rdata = 32'hb7ad8df9;
        1088:    rdata = 32'h854a4595;
        1089:    rdata = 32'h359000ef;
        1090:    rdata = 32'hbf9d4591;
        1091:    rdata = 32'h411cbd61;
        1092:    rdata = 32'hce4e7179;
        1093:    rdata = 32'hd606cc52;
        1094:    rdata = 32'hd226d422;
        1095:    rdata = 32'hca56d04a;
        1096:    rdata = 32'hc65ec85a;
        1097:    rdata = 32'h89b28a2e;
        1098:    rdata = 32'h862eeba5;
        1099:    rdata = 32'h000ef517;
        1100:    rdata = 32'hefc50513;
        1101:    rdata = 32'h26014581;
        1102:    rdata = 32'h000ef517;
        1103:    rdata = 32'hedc50513;
        1104:    rdata = 32'h547000ef;
        1105:    rdata = 32'h000ef417;
        1106:    rdata = 32'hed040413;
        1107:    rdata = 32'h00ef8522;
        1108:    rdata = 32'hdd6d5450;
        1109:    rdata = 32'h1c098413;
        1110:    rdata = 32'h000ef497;
        1111:    rdata = 32'hebc48493;
        1112:    rdata = 32'h85a28526;
        1113:    rdata = 32'h325000ef;
        1114:    rdata = 32'h00ef8526;
        1115:    rdata = 32'h852651d0;
        1116:    rdata = 32'h523000ef;
        1117:    rdata = 32'h0793dd6d;
        1118:    rdata = 32'h9d63fc04;
        1119:    rdata = 32'h50b20089;
        1120:    rdata = 32'h54925422;
        1121:    rdata = 32'h49f25902;
        1122:    rdata = 32'h4ad24a62;
        1123:    rdata = 32'h4bb24b42;
        1124:    rdata = 32'h80826145;
        1125:    rdata = 32'hb7e9843e;
        1126:    rdata = 32'h04134705;
        1127:    rdata = 32'h86631c06;
        1128:    rdata = 32'h4a8506e7;
        1129:    rdata = 32'h02000b13;
        1130:    rdata = 32'h000ef497;
        1131:    rdata = 32'he6c48493;
        1132:    rdata = 32'h493d5bfd;
        1133:    rdata = 32'h012a9633;
        1134:    rdata = 32'h45814781;
        1135:    rdata = 32'h00179693;
        1136:    rdata = 32'hd68396a2;
        1137:    rdata = 32'h97330006;
        1138:    rdata = 32'h8ef100fa;
        1139:    rdata = 32'h8dd9c6dd;
        1140:    rdata = 32'h95e30785;
        1141:    rdata = 32'h8526ff67;
        1142:    rdata = 32'h2ab000ef;
        1143:    rdata = 32'h0a0a1363;
        1144:    rdata = 32'h85264589;
        1145:    rdata = 32'h279000ef;
        1146:    rdata = 32'h8526458d;
        1147:    rdata = 32'h271000ef;
        1148:    rdata = 32'h85264589;
        1149:    rdata = 32'h00ef197d;
        1150:    rdata = 32'h1de32670;
        1151:    rdata = 32'h0793fb79;
        1152:    rdata = 32'h8ee3fc04;
        1153:    rdata = 32'h843ef689;
        1154:    rdata = 32'h862eb76d;
        1155:    rdata = 32'h000ef517;
        1156:    rdata = 32'he1c50513;
        1157:    rdata = 32'h24054585;
        1158:    rdata = 32'h0a934a05;
        1159:    rdata = 32'hf9170200;
        1160:    rdata = 32'h0913000e;
        1161:    rdata = 32'h5b7ddf69;
        1162:    rdata = 32'h163344bd;
        1163:    rdata = 32'h4781009a;
        1164:    rdata = 32'h96934581;
        1165:    rdata = 32'h96a20017;
        1166:    rdata = 32'h0006d683;
        1167:    rdata = 32'h00fa1733;
        1168:    rdata = 32'hca858ef1;
        1169:    rdata = 32'h07858dd9;
        1170:    rdata = 32'hff5795e3;
        1171:    rdata = 32'h00ef854a;
        1172:    rdata = 32'h854a2350;
        1173:    rdata = 32'h43f000ef;
        1174:    rdata = 32'h854add6d;
        1175:    rdata = 32'h00ef14fd;
        1176:    rdata = 32'h94e34290;
        1177:    rdata = 32'h0793fd64;
        1178:    rdata = 32'h8ae3fc04;
        1179:    rdata = 32'h843ef089;
        1180:    rdata = 32'h4713bf65;
        1181:    rdata = 32'h8df9fff7;
        1182:    rdata = 32'h4713b7f9;
        1183:    rdata = 32'h8df9fff7;
        1184:    rdata = 32'h4591bf81;
        1185:    rdata = 32'h00ef8526;
        1186:    rdata = 32'h45951d70;
        1187:    rdata = 32'h00ef8526;
        1188:    rdata = 32'h45911cf0;
        1189:    rdata = 32'hbda5bfb9;
        1190:    rdata = 32'h71397379;
        1191:    rdata = 32'h40030313;
        1192:    rdata = 32'hda26dc22;
        1193:    rdata = 32'hd64ed84a;
        1194:    rdata = 32'hd256d452;
        1195:    rdata = 32'hca66cc62;
        1196:    rdata = 32'hde066a09;
        1197:    rdata = 32'hce5ed05a;
        1198:    rdata = 32'h0818911a;
        1199:    rdata = 32'hc00a0793;
        1200:    rdata = 32'h97ba74fd;
        1201:    rdata = 32'h80048493;
        1202:    rdata = 32'h690994be;
        1203:    rdata = 32'h0613842a;
        1204:    rdata = 32'h45818009;
        1205:    rdata = 32'h10ef8526;
        1206:    rdata = 32'h07930360;
        1207:    rdata = 32'h0818c00a;
        1208:    rdata = 32'h87b397ba;
        1209:    rdata = 32'h7af94127;
        1210:    rdata = 32'hc63e4981;
        1211:    rdata = 32'h60078a13;
        1212:    rdata = 32'h600a8a93;
        1213:    rdata = 32'h60048c13;
        1214:    rdata = 32'h9b134ca1;
        1215:    rdata = 32'h49010109;
        1216:    rdata = 32'h010b5b13;
        1217:    rdata = 32'h4581865a;
        1218:    rdata = 32'h1b938522;
        1219:    rdata = 32'h39590109;
        1220:    rdata = 32'h010bdb93;
        1221:    rdata = 32'h4585865e;
        1222:    rdata = 32'h31698522;
        1223:    rdata = 32'h34798522;
        1224:    rdata = 32'h34898522;
        1225:    rdata = 32'h85a24601;
        1226:    rdata = 32'h34f18552;
        1227:    rdata = 32'h07136709;
        1228:    rdata = 32'h0814c007;
        1229:    rdata = 32'h87a69736;
        1230:    rdata = 32'h86ba9756;
        1231:    rdata = 32'h0c078593;
        1232:    rdata = 32'h0006d603;
        1233:    rdata = 32'h0047d503;
        1234:    rdata = 32'h00c57863;
        1235:    rdata = 32'h01679023;
        1236:    rdata = 32'h01779123;
        1237:    rdata = 32'h00c79223;
        1238:    rdata = 32'h06890799;
        1239:    rdata = 32'hfeb792e3;
        1240:    rdata = 32'h04070713;
        1241:    rdata = 32'hfcfc1be3;
        1242:    rdata = 32'h1de30905;
        1243:    rdata = 32'h0985f999;
        1244:    rdata = 32'hf92995e3;
        1245:    rdata = 32'h07136609;
        1246:    rdata = 32'h0814c006;
        1247:    rdata = 32'h77fd9736;
        1248:    rdata = 32'h059397ba;
        1249:    rdata = 32'h7779c006;
        1250:    rdata = 32'h06130804;
        1251:    rdata = 32'h0513c006;
        1252:    rdata = 32'h95a64007;
        1253:    rdata = 32'h60070713;
        1254:    rdata = 32'h87939626;
        1255:    rdata = 32'h46818027;
        1256:    rdata = 32'h9732952e;
        1257:    rdata = 32'h04000893;
        1258:    rdata = 32'h20000813;
        1259:    rdata = 32'h00d50f33;
        1260:    rdata = 32'h00d70eb3;
        1261:    rdata = 32'h460185be;
        1262:    rdata = 32'hffe5de03;
        1263:    rdata = 32'h00cf0333;
        1264:    rdata = 32'h10230599;
        1265:    rdata = 32'hde0301c3;
        1266:    rdata = 32'h8333ffa5;
        1267:    rdata = 32'h060900ce;
        1268:    rdata = 32'h01c31023;
        1269:    rdata = 32'hff1612e3;
        1270:    rdata = 32'h04068693;
        1271:    rdata = 32'h0c078793;
        1272:    rdata = 32'hfd0696e3;
        1273:    rdata = 32'h08186909;
        1274:    rdata = 32'h079374f9;
        1275:    rdata = 32'h97bac009;
        1276:    rdata = 32'h40048613;
        1277:    rdata = 32'h8522963e;
        1278:    rdata = 32'h3b114581;
        1279:    rdata = 32'h07930818;
        1280:    rdata = 32'h97bac009;
        1281:    rdata = 32'h60048613;
        1282:    rdata = 32'h963e8522;
        1283:    rdata = 32'h33014585;
        1284:    rdata = 32'h3a698522;
        1285:    rdata = 32'h03136309;
        1286:    rdata = 32'h911ac003;
        1287:    rdata = 32'h546250f2;
        1288:    rdata = 32'h594254d2;
        1289:    rdata = 32'h5a2259b2;
        1290:    rdata = 32'h5b025a92;
        1291:    rdata = 32'h4c624bf2;
        1292:    rdata = 32'h61214cd2;
        1293:    rdata = 32'he58d8082;
        1294:    rdata = 32'h0613ee09;
        1295:    rdata = 32'h15970670;
        1296:    rdata = 32'h85930000;
        1297:    rdata = 32'hf5174b25;
        1298:    rdata = 32'h0513000e;
        1299:    rdata = 32'h006fbce5;
        1300:    rdata = 32'h06131810;
        1301:    rdata = 32'h15970670;
        1302:    rdata = 32'h85930000;
        1303:    rdata = 32'hb7e55025;
        1304:    rdata = 32'h9f634785;
        1305:    rdata = 32'he61900f5;
        1306:    rdata = 32'h15974625;
        1307:    rdata = 32'h85930000;
        1308:    rdata = 32'hbfd15565;
        1309:    rdata = 32'h15974625;
        1310:    rdata = 32'h85930000;
        1311:    rdata = 32'hb7e15565;
        1312:    rdata = 32'h46258082;
        1313:    rdata = 32'h00001597;
        1314:    rdata = 32'h55458593;
        1315:    rdata = 32'h000ef517;
        1316:    rdata = 32'hb8850513;
        1317:    rdata = 32'h13b0006f;
        1318:    rdata = 32'h15974625;
        1319:    rdata = 32'h85930000;
        1320:    rdata = 32'hf51754a5;
        1321:    rdata = 32'h0513000e;
        1322:    rdata = 32'h006fb725;
        1323:    rdata = 32'h07131250;
        1324:    rdata = 32'h47830300;
        1325:    rdata = 32'h94630005;
        1326:    rdata = 32'h050500e7;
        1327:    rdata = 32'he391bfdd;
        1328:    rdata = 32'h8082157d;
        1329:    rdata = 32'h00054703;
        1330:    rdata = 32'h02d00793;
        1331:    rdata = 32'h00f71363;
        1332:    rdata = 32'h47250505;
        1333:    rdata = 32'h00054783;
        1334:    rdata = 32'hfd078793;
        1335:    rdata = 32'h0ff7f793;
        1336:    rdata = 32'h00f76863;
        1337:    rdata = 32'h00154783;
        1338:    rdata = 32'hf7ed0505;
        1339:    rdata = 32'h80824505;
        1340:    rdata = 32'h80824501;
        1341:    rdata = 32'h46a50509;
        1342:    rdata = 32'h47834615;
        1343:    rdata = 32'h87130005;
        1344:    rdata = 32'h7713fd07;
        1345:    rdata = 32'hfa630ff7;
        1346:    rdata = 32'hf79300e6;
        1347:    rdata = 32'h8793fdf7;
        1348:    rdata = 32'hf793fbf7;
        1349:    rdata = 32'h68630ff7;
        1350:    rdata = 32'h478300f6;
        1351:    rdata = 32'h05050015;
        1352:    rdata = 32'h4505ffe9;
        1353:    rdata = 32'h45018082;
        1354:    rdata = 32'h87aa8082;
        1355:    rdata = 32'h0005c703;
        1356:    rdata = 32'h07850585;
        1357:    rdata = 32'hfee78fa3;
        1358:    rdata = 32'h8082fb75;
        1359:    rdata = 32'hc68387aa;
        1360:    rdata = 32'h873e0007;
        1361:    rdata = 32'hfee50785;
        1362:    rdata = 32'h0005c783;
        1363:    rdata = 32'h07050585;
        1364:    rdata = 32'hfef70fa3;
        1365:    rdata = 32'h8082fbf5;
        1366:    rdata = 32'h00054783;
        1367:    rdata = 32'h0005c703;
        1368:    rdata = 32'h00e78763;
        1369:    rdata = 32'he963557d;
        1370:    rdata = 32'h450500e7;
        1371:    rdata = 32'hc7818082;
        1372:    rdata = 32'h05850505;
        1373:    rdata = 32'h4501b7d5;
        1374:    rdata = 32'h87aa8082;
        1375:    rdata = 32'h87334501;
        1376:    rdata = 32'h470300a7;
        1377:    rdata = 32'hc3190007;
        1378:    rdata = 32'hbfd50505;
        1379:    rdata = 32'h47898082;
        1380:    rdata = 32'h02f60c63;
        1381:    rdata = 32'h0d634791;
        1382:    rdata = 32'h470502f6;
        1383:    rdata = 32'h14634781;
        1384:    rdata = 32'h079300e6;
        1385:    rdata = 32'h46290640;
        1386:    rdata = 32'hd733cb8d;
        1387:    rdata = 32'h050502f5;
        1388:    rdata = 32'h0ff77693;
        1389:    rdata = 32'h02f686b3;
        1390:    rdata = 32'h03070713;
        1391:    rdata = 32'hfee50fa3;
        1392:    rdata = 32'h02c7d7b3;
        1393:    rdata = 32'hb7cd8d95;
        1394:    rdata = 32'h87936789;
        1395:    rdata = 32'hbfe17107;
        1396:    rdata = 32'h3b9ad7b7;
        1397:    rdata = 32'ha0078793;
        1398:    rdata = 32'h0023b7f9;
        1399:    rdata = 32'h80820005;
        1400:    rdata = 32'hb7754605;
        1401:    rdata = 32'hcc221101;
        1402:    rdata = 32'h842a4611;
        1403:    rdata = 32'hce060048;
        1404:    rdata = 32'h00483f79;
        1405:    rdata = 32'h85aa3d6d;
        1406:    rdata = 32'h3f058522;
        1407:    rdata = 32'h446240f2;
        1408:    rdata = 32'h80826105;
        1409:    rdata = 32'h03000793;
        1410:    rdata = 32'h76130606;
        1411:    rdata = 32'h00230ff6;
        1412:    rdata = 32'h079300f5;
        1413:    rdata = 32'h00a30780;
        1414:    rdata = 32'h482500f5;
        1415:    rdata = 32'hc38587b2;
        1416:    rdata = 32'h00f5f713;
        1417:    rdata = 32'h05770693;
        1418:    rdata = 32'h00e86463;
        1419:    rdata = 32'h03070693;
        1420:    rdata = 32'h00f50733;
        1421:    rdata = 32'h00d700a3;
        1422:    rdata = 32'h17fd8191;
        1423:    rdata = 32'h9532b7cd;
        1424:    rdata = 32'h00050123;
        1425:    rdata = 32'h46058082;
        1426:    rdata = 32'h4611bf75;
        1427:    rdata = 32'h1101bf65;
        1428:    rdata = 32'hce06cc22;
        1429:    rdata = 32'hd563842a;
        1430:    rdata = 32'h07130205;
        1431:    rdata = 32'h002302d0;
        1432:    rdata = 32'h05b300e5;
        1433:    rdata = 32'h461140b0;
        1434:    rdata = 32'h37150048;
        1435:    rdata = 32'h35810048;
        1436:    rdata = 32'h051385aa;
        1437:    rdata = 32'h3d550014;
        1438:    rdata = 32'h446240f2;
        1439:    rdata = 32'h80826105;
        1440:    rdata = 32'h00484611;
        1441:    rdata = 32'h00483729;
        1442:    rdata = 32'h85aa351d;
        1443:    rdata = 32'hb7e58522;
        1444:    rdata = 32'hc4221141;
        1445:    rdata = 32'h842ac606;
        1446:    rdata = 32'he1153535;
        1447:    rdata = 32'h00044703;
        1448:    rdata = 32'h03000793;
        1449:    rdata = 32'h00f71d63;
        1450:    rdata = 32'h00144703;
        1451:    rdata = 32'h07800793;
        1452:    rdata = 32'h00f71763;
        1453:    rdata = 32'h44228522;
        1454:    rdata = 32'h014140b2;
        1455:    rdata = 32'h40b2bd25;
        1456:    rdata = 32'h01414422;
        1457:    rdata = 32'h11418082;
        1458:    rdata = 32'hc606c422;
        1459:    rdata = 32'h3bdd842a;
        1460:    rdata = 32'h00044783;
        1461:    rdata = 32'h0693c91d;
        1462:    rdata = 32'h470102d0;
        1463:    rdata = 32'h00d79463;
        1464:    rdata = 32'h0405872a;
        1465:    rdata = 32'h46294501;
        1466:    rdata = 32'h00044683;
        1467:    rdata = 32'h07b3ca81;
        1468:    rdata = 32'h851302c5;
        1469:    rdata = 32'h0405fd06;
        1470:    rdata = 32'hb7fd953e;
        1471:    rdata = 32'h0533c319;
        1472:    rdata = 32'h40b240a0;
        1473:    rdata = 32'h01414422;
        1474:    rdata = 32'h07138082;
        1475:    rdata = 32'h96630300;
        1476:    rdata = 32'h470304e7;
        1477:    rdata = 32'h07930014;
        1478:    rdata = 32'h10630780;
        1479:    rdata = 32'h852204f7;
        1480:    rdata = 32'hcd053bd1;
        1481:    rdata = 32'h45010409;
        1482:    rdata = 32'h06000713;
        1483:    rdata = 32'h04000693;
        1484:    rdata = 32'h00044783;
        1485:    rdata = 32'h7a63d7f9;
        1486:    rdata = 32'h879300f7;
        1487:    rdata = 32'hf793fa97;
        1488:    rdata = 32'h05120ff7;
        1489:    rdata = 32'h04058d5d;
        1490:    rdata = 32'hf563b7e5;
        1491:    rdata = 32'h879300f6;
        1492:    rdata = 32'hb7f5fc97;
        1493:    rdata = 32'hfd078793;
        1494:    rdata = 32'hc537b7dd;
        1495:    rdata = 32'h0513dead;
        1496:    rdata = 32'hb745eef5;
        1497:    rdata = 32'hfdf57793;
        1498:    rdata = 32'hfbf78793;
        1499:    rdata = 32'h0ff7f793;
        1500:    rdata = 32'h77634765;
        1501:    rdata = 32'h051300f7;
        1502:    rdata = 32'h3513fd05;
        1503:    rdata = 32'h808200a5;
        1504:    rdata = 32'h80824505;
        1505:    rdata = 32'hc4221141;
        1506:    rdata = 32'h06400613;
        1507:    rdata = 32'hf517842a;
        1508:    rdata = 32'h0513000e;
        1509:    rdata = 32'hc6068ae5;
        1510:    rdata = 32'h023000ef;
        1511:    rdata = 32'h852240b2;
        1512:    rdata = 32'h01414422;
        1513:    rdata = 32'h11418082;
        1514:    rdata = 32'h842ac422;
        1515:    rdata = 32'h000ef517;
        1516:    rdata = 32'h89050513;
        1517:    rdata = 32'h00efc606;
        1518:    rdata = 32'h40b20a70;
        1519:    rdata = 32'h44228522;
        1520:    rdata = 32'h80820141;
        1521:    rdata = 32'hc4221141;
        1522:    rdata = 32'hf517842a;
        1523:    rdata = 32'h0513000e;
        1524:    rdata = 32'hc6068725;
        1525:    rdata = 32'h089000ef;
        1526:    rdata = 32'h852240b2;
        1527:    rdata = 32'h01414422;
        1528:    rdata = 32'h418c8082;
        1529:    rdata = 32'hcc221101;
        1530:    rdata = 32'h0048842a;
        1531:    rdata = 32'h3585ce06;
        1532:    rdata = 32'hf517004c;
        1533:    rdata = 32'h0513000e;
        1534:    rdata = 32'h00ef84a5;
        1535:    rdata = 32'h40f20630;
        1536:    rdata = 32'h44628522;
        1537:    rdata = 32'h80826105;
        1538:    rdata = 32'hc4221141;
        1539:    rdata = 32'hf417c606;
        1540:    rdata = 32'h0413000e;
        1541:    rdata = 32'h852282e4;
        1542:    rdata = 32'h003000ef;
        1543:    rdata = 32'h40b2fd6d;
        1544:    rdata = 32'h01414422;
        1545:    rdata = 32'h71758082;
        1546:    rdata = 32'hc326c522;
        1547:    rdata = 32'hdecec14a;
        1548:    rdata = 32'hc706dcd2;
        1549:    rdata = 32'h892e84aa;
        1550:    rdata = 32'h000ef417;
        1551:    rdata = 32'h80440413;
        1552:    rdata = 32'h00001a17;
        1553:    rdata = 32'h7c0a0a13;
        1554:    rdata = 32'h00001997;
        1555:    rdata = 32'h7c498993;
        1556:    rdata = 32'h852285ca;
        1557:    rdata = 32'h009000ef;
        1558:    rdata = 32'h852285d2;
        1559:    rdata = 32'h001000ef;
        1560:    rdata = 32'h8526006c;
        1561:    rdata = 32'h00683705;
        1562:    rdata = 32'he5113525;
        1563:    rdata = 32'h852285ce;
        1564:    rdata = 32'h7ec000ef;
        1565:    rdata = 32'h0068bff1;
        1566:    rdata = 32'h40ba35b9;
        1567:    rdata = 32'h449a442a;
        1568:    rdata = 32'h59f6490a;
        1569:    rdata = 32'h61495a66;
        1570:    rdata = 32'h25738082;
        1571:    rdata = 32'h25f3b000;
        1572:    rdata = 32'h8082b800;
        1573:    rdata = 32'h00010001;
        1574:    rdata = 32'h00010001;
        1575:    rdata = 32'h00010001;
        1576:    rdata = 32'hf9ed15fd;
        1577:    rdata = 32'hc10c8082;
        1578:    rdata = 32'h62f38082;
        1579:    rdata = 32'h80823004;
        1580:    rdata = 32'h300472f3;
        1581:    rdata = 32'hc14c8082;
        1582:    rdata = 32'ha2f362c1;
        1583:    rdata = 32'h80823042;
        1584:    rdata = 32'h00052223;
        1585:    rdata = 32'hb2f362c1;
        1586:    rdata = 32'h80823042;
        1587:    rdata = 32'h02b7c50c;
        1588:    rdata = 32'ha2f30002;
        1589:    rdata = 32'h80823042;
        1590:    rdata = 32'h00052423;
        1591:    rdata = 32'h000202b7;
        1592:    rdata = 32'h3042b2f3;
        1593:    rdata = 32'hc54c8082;
        1594:    rdata = 32'h000402b7;
        1595:    rdata = 32'h3042a2f3;
        1596:    rdata = 32'h26238082;
        1597:    rdata = 32'h02b70005;
        1598:    rdata = 32'hb2f30004;
        1599:    rdata = 32'h80823042;
        1600:    rdata = 32'h02b7c90c;
        1601:    rdata = 32'ha2f30008;
        1602:    rdata = 32'h80823042;
        1603:    rdata = 32'h00052823;
        1604:    rdata = 32'h000802b7;
        1605:    rdata = 32'h3042b2f3;
        1606:    rdata = 32'h71398082;
        1607:    rdata = 32'hde06d036;
        1608:    rdata = 32'hda1adc16;
        1609:    rdata = 32'hd62ad81e;
        1610:    rdata = 32'hd232d42e;
        1611:    rdata = 32'hcc3ece3a;
        1612:    rdata = 32'hc846ca42;
        1613:    rdata = 32'hc476c672;
        1614:    rdata = 32'hc07ec27a;
        1615:    rdata = 32'h000ee697;
        1616:    rdata = 32'h6c46a683;
        1617:    rdata = 32'h2673ce9d;
        1618:    rdata = 32'h42183410;
        1619:    rdata = 32'h8b0d4791;
        1620:    rdata = 32'h4789e311;
        1621:    rdata = 32'h907397b2;
        1622:    rdata = 32'h96823417;
        1623:    rdata = 32'h52e250f2;
        1624:    rdata = 32'h53c25352;
        1625:    rdata = 32'h55a25532;
        1626:    rdata = 32'h56825612;
        1627:    rdata = 32'h47e24772;
        1628:    rdata = 32'h48c24852;
        1629:    rdata = 32'h4ea24e32;
        1630:    rdata = 32'h4f824f12;
        1631:    rdata = 32'h00736121;
        1632:    rdata = 32'ha0013020;
        1633:    rdata = 32'hcc3e7139;
        1634:    rdata = 32'hdc16de06;
        1635:    rdata = 32'hd81eda1a;
        1636:    rdata = 32'hd42ed62a;
        1637:    rdata = 32'hd036d232;
        1638:    rdata = 32'hca42ce3a;
        1639:    rdata = 32'hc672c846;
        1640:    rdata = 32'hc27ac476;
        1641:    rdata = 32'he797c07e;
        1642:    rdata = 32'ha783000e;
        1643:    rdata = 32'h978265e7;
        1644:    rdata = 32'h52e250f2;
        1645:    rdata = 32'h53c25352;
        1646:    rdata = 32'h55a25532;
        1647:    rdata = 32'h56825612;
        1648:    rdata = 32'h47e24772;
        1649:    rdata = 32'h48c24852;
        1650:    rdata = 32'h4ea24e32;
        1651:    rdata = 32'h4f824f12;
        1652:    rdata = 32'h00736121;
        1653:    rdata = 32'h71393020;
        1654:    rdata = 32'hde06cc3e;
        1655:    rdata = 32'hda1adc16;
        1656:    rdata = 32'hd62ad81e;
        1657:    rdata = 32'hd232d42e;
        1658:    rdata = 32'hce3ad036;
        1659:    rdata = 32'hc846ca42;
        1660:    rdata = 32'hc476c672;
        1661:    rdata = 32'hc07ec27a;
        1662:    rdata = 32'h000ee797;
        1663:    rdata = 32'h6107a783;
        1664:    rdata = 32'h50f29782;
        1665:    rdata = 32'h535252e2;
        1666:    rdata = 32'h553253c2;
        1667:    rdata = 32'h561255a2;
        1668:    rdata = 32'h47725682;
        1669:    rdata = 32'h485247e2;
        1670:    rdata = 32'h4e3248c2;
        1671:    rdata = 32'h4f124ea2;
        1672:    rdata = 32'h61214f82;
        1673:    rdata = 32'h30200073;
        1674:    rdata = 32'hcc3e7139;
        1675:    rdata = 32'hdc16de06;
        1676:    rdata = 32'hd81eda1a;
        1677:    rdata = 32'hd42ed62a;
        1678:    rdata = 32'hd036d232;
        1679:    rdata = 32'hca42ce3a;
        1680:    rdata = 32'hc672c846;
        1681:    rdata = 32'hc27ac476;
        1682:    rdata = 32'he797c07e;
        1683:    rdata = 32'ha783000e;
        1684:    rdata = 32'h97825c27;
        1685:    rdata = 32'h52e250f2;
        1686:    rdata = 32'h53c25352;
        1687:    rdata = 32'h55a25532;
        1688:    rdata = 32'h56825612;
        1689:    rdata = 32'h47e24772;
        1690:    rdata = 32'h48c24852;
        1691:    rdata = 32'h4ea24e32;
        1692:    rdata = 32'h4f824f12;
        1693:    rdata = 32'h00736121;
        1694:    rdata = 32'h71393020;
        1695:    rdata = 32'hde06cc3e;
        1696:    rdata = 32'hda1adc16;
        1697:    rdata = 32'hd62ad81e;
        1698:    rdata = 32'hd232d42e;
        1699:    rdata = 32'hce3ad036;
        1700:    rdata = 32'hc846ca42;
        1701:    rdata = 32'hc476c672;
        1702:    rdata = 32'hc07ec27a;
        1703:    rdata = 32'h000ee797;
        1704:    rdata = 32'h5747a783;
        1705:    rdata = 32'h50f29782;
        1706:    rdata = 32'h535252e2;
        1707:    rdata = 32'h553253c2;
        1708:    rdata = 32'h561255a2;
        1709:    rdata = 32'h47725682;
        1710:    rdata = 32'h485247e2;
        1711:    rdata = 32'h4e3248c2;
        1712:    rdata = 32'h4f124ea2;
        1713:    rdata = 32'h61214f82;
        1714:    rdata = 32'h30200073;
        1715:    rdata = 32'h8082c10c;
        1716:    rdata = 32'h00163613;
        1717:    rdata = 32'h000ee517;
        1718:    rdata = 32'h56050513;
        1719:    rdata = 32'h1141a8e9;
        1720:    rdata = 32'h000ee517;
        1721:    rdata = 32'h55450513;
        1722:    rdata = 32'h28c5c606;
        1723:    rdata = 32'h157d40b2;
        1724:    rdata = 32'h00a03533;
        1725:    rdata = 32'h80820141;
        1726:    rdata = 32'h87324108;
        1727:    rdata = 32'h862e4685;
        1728:    rdata = 32'h006f4581;
        1729:    rdata = 32'h11016480;
        1730:    rdata = 32'hc62ecc22;
        1731:    rdata = 32'hce06842a;
        1732:    rdata = 32'h87aa37f9;
        1733:    rdata = 32'h40084632;
        1734:    rdata = 32'h45814685;
        1735:    rdata = 32'h4591c391;
        1736:    rdata = 32'h40f22d29;
        1737:    rdata = 32'h35334462;
        1738:    rdata = 32'h610500a0;
        1739:    rdata = 32'h41088082;
        1740:    rdata = 32'h4685862e;
        1741:    rdata = 32'h006f4581;
        1742:    rdata = 32'h41086300;
        1743:    rdata = 32'h4705862e;
        1744:    rdata = 32'h45a14685;
        1745:    rdata = 32'h4108a519;
        1746:    rdata = 32'h4701862e;
        1747:    rdata = 32'h45a14685;
        1748:    rdata = 32'h4108abed;
        1749:    rdata = 32'h862e1141;
        1750:    rdata = 32'h45b14685;
        1751:    rdata = 32'h2bf1c606;
        1752:    rdata = 32'h353340b2;
        1753:    rdata = 32'h014100a0;
        1754:    rdata = 32'h41088082;
        1755:    rdata = 32'h4701862e;
        1756:    rdata = 32'h45b14685;
        1757:    rdata = 32'h4108abd9;
        1758:    rdata = 32'h4705862e;
        1759:    rdata = 32'h45c14685;
        1760:    rdata = 32'h4108a3e9;
        1761:    rdata = 32'h4701862e;
        1762:    rdata = 32'h45c14685;
        1763:    rdata = 32'h4108ab7d;
        1764:    rdata = 32'h862e1141;
        1765:    rdata = 32'h45d14685;
        1766:    rdata = 32'h2345c606;
        1767:    rdata = 32'h353340b2;
        1768:    rdata = 32'h014100a0;
        1769:    rdata = 32'h41088082;
        1770:    rdata = 32'h4701862e;
        1771:    rdata = 32'h45d14685;
        1772:    rdata = 32'hc10cab69;
        1773:    rdata = 32'h47bd8082;
        1774:    rdata = 32'h87324108;
        1775:    rdata = 32'h00b7e863;
        1776:    rdata = 32'hf6130586;
        1777:    rdata = 32'h468d0fe5;
        1778:    rdata = 32'ha3414581;
        1779:    rdata = 32'h058615c1;
        1780:    rdata = 32'h0fe5f613;
        1781:    rdata = 32'h4591468d;
        1782:    rdata = 32'h1141bfcd;
        1783:    rdata = 32'h47bdc606;
        1784:    rdata = 32'he6634108;
        1785:    rdata = 32'h961302b7;
        1786:    rdata = 32'h468d0015;
        1787:    rdata = 32'h0fe67613;
        1788:    rdata = 32'h23a14581;
        1789:    rdata = 32'h470587aa;
        1790:    rdata = 32'h87634505;
        1791:    rdata = 32'h470900e7;
        1792:    rdata = 32'h93634501;
        1793:    rdata = 32'h450900e7;
        1794:    rdata = 32'h014140b2;
        1795:    rdata = 32'h86138082;
        1796:    rdata = 32'h0606ff05;
        1797:    rdata = 32'h7613468d;
        1798:    rdata = 32'h45910fe6;
        1799:    rdata = 32'h6785bfd9;
        1800:    rdata = 32'h0613c10c;
        1801:    rdata = 32'h95be4000;
        1802:    rdata = 32'ha1fd0511;
        1803:    rdata = 32'h872e4108;
        1804:    rdata = 32'h46094685;
        1805:    rdata = 32'hab114581;
        1806:    rdata = 32'h872e4108;
        1807:    rdata = 32'h460d4685;
        1808:    rdata = 32'ha3214581;
        1809:    rdata = 32'h872e4108;
        1810:    rdata = 32'h46114685;
        1811:    rdata = 32'ha9f54581;
        1812:    rdata = 32'h872e4108;
        1813:    rdata = 32'h46154685;
        1814:    rdata = 32'ha9c54581;
        1815:    rdata = 32'hc78c411c;
        1816:    rdata = 32'h411c8082;
        1817:    rdata = 32'h808247c8;
        1818:    rdata = 32'h11414108;
        1819:    rdata = 32'h0ff00693;
        1820:    rdata = 32'h45914605;
        1821:    rdata = 32'h21d1c606;
        1822:    rdata = 32'h751340b2;
        1823:    rdata = 32'h01410ff5;
        1824:    rdata = 32'h411c8082;
        1825:    rdata = 32'h8082cb8c;
        1826:    rdata = 32'h06134108;
        1827:    rdata = 32'h05410400;
        1828:    rdata = 32'h411ca385;
        1829:    rdata = 32'h80824ba8;
        1830:    rdata = 32'h410c87ae;
        1831:    rdata = 32'h04000613;
        1832:    rdata = 32'h8593853e;
        1833:    rdata = 32'ha3a90505;
        1834:    rdata = 32'h872e4108;
        1835:    rdata = 32'h03f00693;
        1836:    rdata = 32'h05934601;
        1837:    rdata = 32'ha9511000;
        1838:    rdata = 32'h872e4108;
        1839:    rdata = 32'h03f00693;
        1840:    rdata = 32'h05934619;
        1841:    rdata = 32'ha1511000;
        1842:    rdata = 32'h872e4108;
        1843:    rdata = 32'h07f00693;
        1844:    rdata = 32'h05934601;
        1845:    rdata = 32'ha9951080;
        1846:    rdata = 32'h872e4108;
        1847:    rdata = 32'h03f00693;
        1848:    rdata = 32'h05934631;
        1849:    rdata = 32'ha1951000;
        1850:    rdata = 32'h872e4108;
        1851:    rdata = 32'h03f00693;
        1852:    rdata = 32'h05934649;
        1853:    rdata = 32'ha9911000;
        1854:    rdata = 32'h872e4108;
        1855:    rdata = 32'h03f00693;
        1856:    rdata = 32'h05934661;
        1857:    rdata = 32'ha1911000;
        1858:    rdata = 32'h872e4108;
        1859:    rdata = 32'h03f00693;
        1860:    rdata = 32'h05934601;
        1861:    rdata = 32'ha9151040;
        1862:    rdata = 32'h872e4108;
        1863:    rdata = 32'h03f00693;
        1864:    rdata = 32'h05934619;
        1865:    rdata = 32'ha1151040;
        1866:    rdata = 32'h872e4108;
        1867:    rdata = 32'h03f00693;
        1868:    rdata = 32'h05934631;
        1869:    rdata = 32'ha9111040;
        1870:    rdata = 32'h872e4108;
        1871:    rdata = 32'h03f00693;
        1872:    rdata = 32'h05934649;
        1873:    rdata = 32'ha1111040;
        1874:    rdata = 32'h872e4108;
        1875:    rdata = 32'h03f00693;
        1876:    rdata = 32'h05934661;
        1877:    rdata = 32'haed51040;
        1878:    rdata = 32'h872e4108;
        1879:    rdata = 32'h0ff00693;
        1880:    rdata = 32'h05934639;
        1881:    rdata = 32'ha6d51080;
        1882:    rdata = 32'h872e4108;
        1883:    rdata = 32'h0ff00693;
        1884:    rdata = 32'h05934659;
        1885:    rdata = 32'haed11080;
        1886:    rdata = 32'h872e4108;
        1887:    rdata = 32'h07f00693;
        1888:    rdata = 32'h0593461d;
        1889:    rdata = 32'ha6d11080;
        1890:    rdata = 32'h872e4108;
        1891:    rdata = 32'h46094685;
        1892:    rdata = 32'h20000593;
        1893:    rdata = 32'h4108ae5d;
        1894:    rdata = 32'h4685872e;
        1895:    rdata = 32'h05934605;
        1896:    rdata = 32'ha6652000;
        1897:    rdata = 32'h872e4108;
        1898:    rdata = 32'h460d469d;
        1899:    rdata = 32'h20000593;
        1900:    rdata = 32'h4108ae69;
        1901:    rdata = 32'h4685872e;
        1902:    rdata = 32'h05934601;
        1903:    rdata = 32'ha6712000;
        1904:    rdata = 32'hc7134108;
        1905:    rdata = 32'h46850015;
        1906:    rdata = 32'h45814601;
        1907:    rdata = 32'h7139aebd;
        1908:    rdata = 32'h89aed64e;
        1909:    rdata = 32'hdc224585;
        1910:    rdata = 32'hd84ada26;
        1911:    rdata = 32'hd256d452;
        1912:    rdata = 32'hce5ed05a;
        1913:    rdata = 32'h893284aa;
        1914:    rdata = 32'h3fd9de06;
        1915:    rdata = 32'h44334791;
        1916:    rdata = 32'h4a0102f9;
        1917:    rdata = 32'h4b914a81;
        1918:    rdata = 32'h00448b13;
        1919:    rdata = 32'h028ad763;
        1920:    rdata = 32'h86334781;
        1921:    rdata = 32'h06b30149;
        1922:    rdata = 32'hc68300f6;
        1923:    rdata = 32'h00780006;
        1924:    rdata = 32'h0023973e;
        1925:    rdata = 32'h078500d7;
        1926:    rdata = 32'hff7797e3;
        1927:    rdata = 32'h85d24632;
        1928:    rdata = 32'h2621855a;
        1929:    rdata = 32'h0a110a85;
        1930:    rdata = 32'h87a2bfd1;
        1931:    rdata = 32'h00045363;
        1932:    rdata = 32'h95934781;
        1933:    rdata = 32'h05330027;
        1934:    rdata = 32'h096340b9;
        1935:    rdata = 32'h478102b9;
        1936:    rdata = 32'h4701468d;
        1937:    rdata = 32'h00a7d763;
        1938:    rdata = 32'h00f58733;
        1939:    rdata = 32'h4703974e;
        1940:    rdata = 32'h00700007;
        1941:    rdata = 32'h0023963e;
        1942:    rdata = 32'h078500e6;
        1943:    rdata = 32'hfed793e3;
        1944:    rdata = 32'h000107a3;
        1945:    rdata = 32'h85134632;
        1946:    rdata = 32'h24c10044;
        1947:    rdata = 32'h50f25462;
        1948:    rdata = 32'h59b25942;
        1949:    rdata = 32'h5a925a22;
        1950:    rdata = 32'h4bf25b02;
        1951:    rdata = 32'h54d28526;
        1952:    rdata = 32'h61214581;
        1953:    rdata = 32'h4108bf35;
        1954:    rdata = 32'h46854705;
        1955:    rdata = 32'h45814605;
        1956:    rdata = 32'h4108ac6d;
        1957:    rdata = 32'h46851141;
        1958:    rdata = 32'h45914601;
        1959:    rdata = 32'h2c71c606;
        1960:    rdata = 32'h353340b2;
        1961:    rdata = 32'h014100a0;
        1962:    rdata = 32'hc10c8082;
        1963:    rdata = 32'h411c8082;
        1964:    rdata = 32'h8082c7cc;
        1965:    rdata = 32'h47054108;
        1966:    rdata = 32'h46014685;
        1967:    rdata = 32'ha4714581;
        1968:    rdata = 32'h47014108;
        1969:    rdata = 32'h46014685;
        1970:    rdata = 32'ha4414581;
        1971:    rdata = 32'h47014108;
        1972:    rdata = 32'h46014685;
        1973:    rdata = 32'hac954591;
        1974:    rdata = 32'h47014108;
        1975:    rdata = 32'h46014685;
        1976:    rdata = 32'ha4a545c1;
        1977:    rdata = 32'h11414108;
        1978:    rdata = 32'h46014685;
        1979:    rdata = 32'hc60645d1;
        1980:    rdata = 32'h40b224a9;
        1981:    rdata = 32'h00a03533;
        1982:    rdata = 32'h80820141;
        1983:    rdata = 32'h47014108;
        1984:    rdata = 32'h46014685;
        1985:    rdata = 32'ha49145d1;
        1986:    rdata = 32'hc4221141;
        1987:    rdata = 32'h842ac606;
        1988:    rdata = 32'h400837f5;
        1989:    rdata = 32'h40b24422;
        1990:    rdata = 32'h46854705;
        1991:    rdata = 32'h45c14601;
        1992:    rdata = 32'ha4250141;
        1993:    rdata = 32'h8082c10c;
        1994:    rdata = 32'hc4221141;
        1995:    rdata = 32'h4108842a;
        1996:    rdata = 32'h06934731;
        1997:    rdata = 32'h46010ff0;
        1998:    rdata = 32'hc60645c1;
        1999:    rdata = 32'h46092439;
        2000:    rdata = 32'he51745fd;
        2001:    rdata = 32'h0513000e;
        2002:    rdata = 32'hf0ef0f25;
        2003:    rdata = 32'h4609c6df;
        2004:    rdata = 32'he51745f9;
        2005:    rdata = 32'h0513000e;
        2006:    rdata = 32'hf0ef0e25;
        2007:    rdata = 32'h4008c5df;
        2008:    rdata = 32'h40b24422;
        2009:    rdata = 32'h46854705;
        2010:    rdata = 32'h45814601;
        2011:    rdata = 32'haaf10141;
        2012:    rdata = 32'h11414108;
        2013:    rdata = 32'h46014685;
        2014:    rdata = 32'hc6064591;
        2015:    rdata = 32'h40b22a7d;
        2016:    rdata = 32'h00a03533;
        2017:    rdata = 32'h80820141;
        2018:    rdata = 32'h11414108;
        2019:    rdata = 32'h0ff00693;
        2020:    rdata = 32'h45b14601;
        2021:    rdata = 32'h2255c606;
        2022:    rdata = 32'h751340b2;
        2023:    rdata = 32'h01410ff5;
        2024:    rdata = 32'h11418082;
        2025:    rdata = 32'hc606c422;
        2026:    rdata = 32'h8522842a;
        2027:    rdata = 32'hdd7537d1;
        2028:    rdata = 32'h44228522;
        2029:    rdata = 32'h014140b2;
        2030:    rdata = 32'h1101bfc1;
        2031:    rdata = 32'hca26cc22;
        2032:    rdata = 32'hc64ec84a;
        2033:    rdata = 32'hc05ac256;
        2034:    rdata = 32'hc452ce06;
        2035:    rdata = 32'h892e84aa;
        2036:    rdata = 32'h440189b2;
        2037:    rdata = 32'h4b214aa9;
        2038:    rdata = 32'h03345f63;
        2039:    rdata = 32'h0a338526;
        2040:    rdata = 32'h37c10089;
        2041:    rdata = 32'h00aa0023;
        2042:    rdata = 32'h01551f63;
        2043:    rdata = 32'h000a0023;
        2044:    rdata = 32'h40f24501;
        2045:    rdata = 32'h44d24462;
        2046:    rdata = 32'h49b24942;
        2047:    rdata = 32'h4a924a22;
        2048:    rdata = 32'h61054b02;
        2049:    rdata = 32'h14638082;
        2050:    rdata = 32'hc4010165;
        2051:    rdata = 32'h04051479;
        2052:    rdata = 32'h547db7e1;
        2053:    rdata = 32'h4505bfed;
        2054:    rdata = 32'h4108bfe9;
        2055:    rdata = 32'h46851141;
        2056:    rdata = 32'h45914605;
        2057:    rdata = 32'h2a11c606;
        2058:    rdata = 32'h353340b2;
        2059:    rdata = 32'h014100a0;
        2060:    rdata = 32'h41088082;
        2061:    rdata = 32'h0693872e;
        2062:    rdata = 32'h46010ff0;
        2063:    rdata = 32'ha23145a1;
        2064:    rdata = 32'hcc221101;
        2065:    rdata = 32'h842ace06;
        2066:    rdata = 32'hc62e8522;
        2067:    rdata = 32'h45b237f9;
        2068:    rdata = 32'h8522fd65;
        2069:    rdata = 32'h40f24462;
        2070:    rdata = 32'hbfe16105;
        2071:    rdata = 32'hc4221141;
        2072:    rdata = 32'hc606c226;
        2073:    rdata = 32'h842e84aa;
        2074:    rdata = 32'h00044583;
        2075:    rdata = 32'h8526c589;
        2076:    rdata = 32'h37f90405;
        2077:    rdata = 32'h40b2bfd5;
        2078:    rdata = 32'h44924422;
        2079:    rdata = 32'h80820141;
        2080:    rdata = 32'h47014108;
        2081:    rdata = 32'h46014685;
        2082:    rdata = 32'ha0c145d1;
        2083:    rdata = 32'h11414108;
        2084:    rdata = 32'h46014685;
        2085:    rdata = 32'hc60645e1;
        2086:    rdata = 32'h40b2204d;
        2087:    rdata = 32'h00a03533;
        2088:    rdata = 32'h80820141;
        2089:    rdata = 32'h47014108;
        2090:    rdata = 32'h46014685;
        2091:    rdata = 32'ha87145e1;
        2092:    rdata = 32'hc4221141;
        2093:    rdata = 32'h842ac606;
        2094:    rdata = 32'h400837f5;
        2095:    rdata = 32'h40b24422;
        2096:    rdata = 32'h46854705;
        2097:    rdata = 32'h45d14601;
        2098:    rdata = 32'ha0410141;
        2099:    rdata = 32'h47014108;
        2100:    rdata = 32'h46054685;
        2101:    rdata = 32'ha89545d1;
        2102:    rdata = 32'h11414108;
        2103:    rdata = 32'h46054685;
        2104:    rdata = 32'hc60645e1;
        2105:    rdata = 32'h40b22899;
        2106:    rdata = 32'h00a03533;
        2107:    rdata = 32'h80820141;
        2108:    rdata = 32'h47014108;
        2109:    rdata = 32'h46054685;
        2110:    rdata = 32'ha88145e1;
        2111:    rdata = 32'hc4221141;
        2112:    rdata = 32'h842ac606;
        2113:    rdata = 32'h400837f5;
        2114:    rdata = 32'h40b24422;
        2115:    rdata = 32'h46854705;
        2116:    rdata = 32'h45d14605;
        2117:    rdata = 32'ha8150141;
        2118:    rdata = 32'hc150c10c;
        2119:    rdata = 32'hf7938082;
        2120:    rdata = 32'h410cffc5;
        2121:    rdata = 32'h418895be;
        2122:    rdata = 32'hf7938082;
        2123:    rdata = 32'h410cffc5;
        2124:    rdata = 32'hc19095be;
        2125:    rdata = 32'h41488082;
        2126:    rdata = 32'h99f18082;
        2127:    rdata = 32'h411c952e;
        2128:    rdata = 32'h00c7d7b3;
        2129:    rdata = 32'h00d7f533;
        2130:    rdata = 32'h99f18082;
        2131:    rdata = 32'h410c952e;
        2132:    rdata = 32'h00c697b3;
        2133:    rdata = 32'hfff7c793;
        2134:    rdata = 32'h8fed8ef9;
        2135:    rdata = 32'h00c696b3;
        2136:    rdata = 32'hc1148edd;
        2137:    rdata = 32'h99f18082;
        2138:    rdata = 32'h411c952e;
        2139:    rdata = 32'h00c696b3;
        2140:    rdata = 32'hc1148ebd;
        2141:    rdata = 32'h00008082;
        2142:    rdata = 32'h00300793;
        2143:    rdata = 32'h02c7f863;
        2144:    rdata = 32'h00b567b3;
        2145:    rdata = 32'h0037f793;
        2146:    rdata = 32'h00300693;
        2147:    rdata = 32'h04079e63;
        2148:    rdata = 32'h00052703;
        2149:    rdata = 32'h0005a783;
        2150:    rdata = 32'h04f71863;
        2151:    rdata = 32'hffc60613;
        2152:    rdata = 32'h00450513;
        2153:    rdata = 32'h00458593;
        2154:    rdata = 32'hfec6e4e3;
        2155:    rdata = 32'hfff60693;
        2156:    rdata = 32'h02060863;
        2157:    rdata = 32'h00168693;
        2158:    rdata = 32'h00d506b3;
        2159:    rdata = 32'h0080006f;
        2160:    rdata = 32'h02d50063;
        2161:    rdata = 32'h00054783;
        2162:    rdata = 32'h0005c703;
        2163:    rdata = 32'h00150513;
        2164:    rdata = 32'h00158593;
        2165:    rdata = 32'hfee786e3;
        2166:    rdata = 32'h40e78533;
        2167:    rdata = 32'h00008067;
        2168:    rdata = 32'h00000513;
        2169:    rdata = 32'h00008067;
        2170:    rdata = 32'hfff60693;
        2171:    rdata = 32'hfc9ff06f;
        2172:    rdata = 32'h00a5c7b3;
        2173:    rdata = 32'h0037f793;
        2174:    rdata = 32'h00c508b3;
        2175:    rdata = 32'h06079263;
        2176:    rdata = 32'h00300793;
        2177:    rdata = 32'h04c7fe63;
        2178:    rdata = 32'h00357793;
        2179:    rdata = 32'h00050713;
        2180:    rdata = 32'h06079863;
        2181:    rdata = 32'hffc8f613;
        2182:    rdata = 32'hfe060793;
        2183:    rdata = 32'h08f76c63;
        2184:    rdata = 32'h02c77c63;
        2185:    rdata = 32'h00058693;
        2186:    rdata = 32'h00070793;
        2187:    rdata = 32'h0006a803;
        2188:    rdata = 32'h00478793;
        2189:    rdata = 32'h00468693;
        2190:    rdata = 32'hff07ae23;
        2191:    rdata = 32'hfec7e8e3;
        2192:    rdata = 32'hfff60793;
        2193:    rdata = 32'h40e787b3;
        2194:    rdata = 32'hffc7f793;
        2195:    rdata = 32'h00478793;
        2196:    rdata = 32'h00f70733;
        2197:    rdata = 32'h00f585b3;
        2198:    rdata = 32'h01176863;
        2199:    rdata = 32'h00008067;
        2200:    rdata = 32'h00050713;
        2201:    rdata = 32'hff157ce3;
        2202:    rdata = 32'h0005c783;
        2203:    rdata = 32'h00170713;
        2204:    rdata = 32'h00158593;
        2205:    rdata = 32'hfef70fa3;
        2206:    rdata = 32'hff1768e3;
        2207:    rdata = 32'h00008067;
        2208:    rdata = 32'h0005c683;
        2209:    rdata = 32'h00170713;
        2210:    rdata = 32'h00377793;
        2211:    rdata = 32'hfed70fa3;
        2212:    rdata = 32'h00158593;
        2213:    rdata = 32'hf80780e3;
        2214:    rdata = 32'h0005c683;
        2215:    rdata = 32'h00170713;
        2216:    rdata = 32'h00377793;
        2217:    rdata = 32'hfed70fa3;
        2218:    rdata = 32'h00158593;
        2219:    rdata = 32'hfc079ae3;
        2220:    rdata = 32'hf65ff06f;
        2221:    rdata = 32'h0045a683;
        2222:    rdata = 32'h0005a283;
        2223:    rdata = 32'h0085af83;
        2224:    rdata = 32'h00c5af03;
        2225:    rdata = 32'h0105ae83;
        2226:    rdata = 32'h0145ae03;
        2227:    rdata = 32'h0185a303;
        2228:    rdata = 32'h01c5a803;
        2229:    rdata = 32'h00d72223;
        2230:    rdata = 32'h0205a683;
        2231:    rdata = 32'h00572023;
        2232:    rdata = 32'h01f72423;
        2233:    rdata = 32'h01e72623;
        2234:    rdata = 32'h01d72823;
        2235:    rdata = 32'h01c72a23;
        2236:    rdata = 32'h00672c23;
        2237:    rdata = 32'h01072e23;
        2238:    rdata = 32'h02d72023;
        2239:    rdata = 32'h02470713;
        2240:    rdata = 32'h02458593;
        2241:    rdata = 32'hfaf768e3;
        2242:    rdata = 32'hf19ff06f;
        2243:    rdata = 32'h00f00313;
        2244:    rdata = 32'h00050713;
        2245:    rdata = 32'h02c37e63;
        2246:    rdata = 32'h00f77793;
        2247:    rdata = 32'h0a079063;
        2248:    rdata = 32'h08059263;
        2249:    rdata = 32'hff067693;
        2250:    rdata = 32'h00f67613;
        2251:    rdata = 32'h00e686b3;
        2252:    rdata = 32'h00b72023;
        2253:    rdata = 32'h00b72223;
        2254:    rdata = 32'h00b72423;
        2255:    rdata = 32'h00b72623;
        2256:    rdata = 32'h01070713;
        2257:    rdata = 32'hfed766e3;
        2258:    rdata = 32'h00061463;
        2259:    rdata = 32'h00008067;
        2260:    rdata = 32'h40c306b3;
        2261:    rdata = 32'h00269693;
        2262:    rdata = 32'h00000297;
        2263:    rdata = 32'h005686b3;
        2264:    rdata = 32'h00c68067;
        2265:    rdata = 32'h00b70723;
        2266:    rdata = 32'h00b706a3;
        2267:    rdata = 32'h00b70623;
        2268:    rdata = 32'h00b705a3;
        2269:    rdata = 32'h00b70523;
        2270:    rdata = 32'h00b704a3;
        2271:    rdata = 32'h00b70423;
        2272:    rdata = 32'h00b703a3;
        2273:    rdata = 32'h00b70323;
        2274:    rdata = 32'h00b702a3;
        2275:    rdata = 32'h00b70223;
        2276:    rdata = 32'h00b701a3;
        2277:    rdata = 32'h00b70123;
        2278:    rdata = 32'h00b700a3;
        2279:    rdata = 32'h00b70023;
        2280:    rdata = 32'h00008067;
        2281:    rdata = 32'h0ff5f593;
        2282:    rdata = 32'h00859693;
        2283:    rdata = 32'h00d5e5b3;
        2284:    rdata = 32'h01059693;
        2285:    rdata = 32'h00d5e5b3;
        2286:    rdata = 32'hf6dff06f;
        2287:    rdata = 32'h00279693;
        2288:    rdata = 32'h00000297;
        2289:    rdata = 32'h005686b3;
        2290:    rdata = 32'h00008293;
        2291:    rdata = 32'hfa0680e7;
        2292:    rdata = 32'h00028093;
        2293:    rdata = 32'hff078793;
        2294:    rdata = 32'h40f70733;
        2295:    rdata = 32'h00f60633;
        2296:    rdata = 32'hf6c378e3;
        2297:    rdata = 32'hf3dff06f;
        2298:    rdata = 32'hc4221141;
        2299:    rdata = 32'hc04ac226;
        2300:    rdata = 32'h842ac606;
        2301:    rdata = 32'h84b2892e;
        2302:    rdata = 32'h01240e63;
        2303:    rdata = 32'h04000613;
        2304:    rdata = 32'h852285a6;
        2305:    rdata = 32'hd75ff0ef;
        2306:    rdata = 32'h0413ed09;
        2307:    rdata = 32'h84930404;
        2308:    rdata = 32'hb7dd0404;
        2309:    rdata = 32'h40b24505;
        2310:    rdata = 32'h44924422;
        2311:    rdata = 32'h01414902;
        2312:    rdata = 32'h45018082;
        2313:    rdata = 32'h1101bfcd;
        2314:    rdata = 32'h00001597;
        2315:    rdata = 32'hbb858593;
        2316:    rdata = 32'h000ee517;
        2317:    rdata = 32'hbfc50513;
        2318:    rdata = 32'hf0efce06;
        2319:    rdata = 32'h0068b8af;
        2320:    rdata = 32'hb74fe0ef;
        2321:    rdata = 32'h450140f2;
        2322:    rdata = 32'h80826105;
        2323:    rdata = 32'h010017b7;
        2324:    rdata = 32'h000ee717;
        2325:    rdata = 32'hbef72023;
        2326:    rdata = 32'h07b78082;
        2327:    rdata = 32'he7170100;
        2328:    rdata = 32'h2b23000e;
        2329:    rdata = 32'h8082bcf7;
        2330:    rdata = 32'h010105b7;
        2331:    rdata = 32'h000ee517;
        2332:    rdata = 32'hba850513;
        2333:    rdata = 32'hfaaff06f;
        2334:    rdata = 32'h010047b7;
        2335:    rdata = 32'h000ee717;
        2336:    rdata = 32'hbaf72e23;
        2337:    rdata = 32'h27b78082;
        2338:    rdata = 32'he7170100;
        2339:    rdata = 32'h2923000e;
        2340:    rdata = 32'h8082baf7;
        2341:    rdata = 32'h00000000;
        2342:    rdata = 32'h00000000;
        2343:    rdata = 32'h00000000;
        2344:    rdata = 32'h00000000;
        2345:    rdata = 32'h0001244c;
        2346:    rdata = 32'h0001245a;
        2347:    rdata = 32'h00012468;
        2348:    rdata = 32'h00012478;
        2349:    rdata = 32'h00012486;
        2350:    rdata = 32'hffffe372;
        2351:    rdata = 32'hffffe378;
        2352:    rdata = 32'hffffe37e;
        2353:    rdata = 32'hffffe384;
        2354:    rdata = 32'hffffe392;
        2355:    rdata = 32'hffffe39a;
        2356:    rdata = 32'hffffe3a2;
        2357:    rdata = 32'hffffe3aa;
        2358:    rdata = 32'hffffe3b2;
        2359:    rdata = 32'hffffe3ba;
        2360:    rdata = 32'hffffe3c2;
        2361:    rdata = 32'hffffe3c8;
        2362:    rdata = 32'hffffe3ce;
        2363:    rdata = 32'hffffe3d4;
        2364:    rdata = 32'h00010000;
        2365:    rdata = 32'h00030002;
        2366:    rdata = 32'h00050004;
        2367:    rdata = 32'h00070006;
        2368:    rdata = 32'h00090008;
        2369:    rdata = 32'h000b000a;
        2370:    rdata = 32'h000d000c;
        2371:    rdata = 32'h000f000e;
        2372:    rdata = 32'h00110010;
        2373:    rdata = 32'h00130012;
        2374:    rdata = 32'h00150014;
        2375:    rdata = 32'h00170016;
        2376:    rdata = 32'h00190018;
        2377:    rdata = 32'h001b001a;
        2378:    rdata = 32'h001d001c;
        2379:    rdata = 32'h001f001e;
        2380:    rdata = 32'h00210020;
        2381:    rdata = 32'h00230022;
        2382:    rdata = 32'h00250024;
        2383:    rdata = 32'h00270026;
        2384:    rdata = 32'h00290028;
        2385:    rdata = 32'h002b002a;
        2386:    rdata = 32'h002d002c;
        2387:    rdata = 32'h002f002e;
        2388:    rdata = 32'h00310030;
        2389:    rdata = 32'h00330032;
        2390:    rdata = 32'h00350034;
        2391:    rdata = 32'h00370036;
        2392:    rdata = 32'h00390038;
        2393:    rdata = 32'h003b003a;
        2394:    rdata = 32'h003d003c;
        2395:    rdata = 32'h003f003e;
        2396:    rdata = 32'h00410040;
        2397:    rdata = 32'h00430042;
        2398:    rdata = 32'h00450044;
        2399:    rdata = 32'h00470046;
        2400:    rdata = 32'h00490048;
        2401:    rdata = 32'h004b004a;
        2402:    rdata = 32'h004d004c;
        2403:    rdata = 32'h004f004e;
        2404:    rdata = 32'h00510050;
        2405:    rdata = 32'h00530052;
        2406:    rdata = 32'h00550054;
        2407:    rdata = 32'h00570056;
        2408:    rdata = 32'h00590058;
        2409:    rdata = 32'h005b005a;
        2410:    rdata = 32'h005d005c;
        2411:    rdata = 32'h005f005e;
        2412:    rdata = 32'h00610060;
        2413:    rdata = 32'h00630062;
        2414:    rdata = 32'h00650064;
        2415:    rdata = 32'h00670066;
        2416:    rdata = 32'h00690068;
        2417:    rdata = 32'h006b006a;
        2418:    rdata = 32'h006d006c;
        2419:    rdata = 32'h006f006e;
        2420:    rdata = 32'h00710070;
        2421:    rdata = 32'h00730072;
        2422:    rdata = 32'h00750074;
        2423:    rdata = 32'h00770076;
        2424:    rdata = 32'h00790078;
        2425:    rdata = 32'h007b007a;
        2426:    rdata = 32'h007d007c;
        2427:    rdata = 32'h007f007e;
        2428:    rdata = 32'h00810080;
        2429:    rdata = 32'h00830082;
        2430:    rdata = 32'h00850084;
        2431:    rdata = 32'h00870086;
        2432:    rdata = 32'h00890088;
        2433:    rdata = 32'h008b008a;
        2434:    rdata = 32'h008d008c;
        2435:    rdata = 32'h008f008e;
        2436:    rdata = 32'h00910090;
        2437:    rdata = 32'h00930092;
        2438:    rdata = 32'h00950094;
        2439:    rdata = 32'h00970096;
        2440:    rdata = 32'h00990098;
        2441:    rdata = 32'h009b009a;
        2442:    rdata = 32'h009d009c;
        2443:    rdata = 32'h009f009e;
        2444:    rdata = 32'h00a100a0;
        2445:    rdata = 32'h00a300a2;
        2446:    rdata = 32'h00a500a4;
        2447:    rdata = 32'h00a700a6;
        2448:    rdata = 32'h00a900a8;
        2449:    rdata = 32'h00ab00aa;
        2450:    rdata = 32'h00ad00ac;
        2451:    rdata = 32'h00af00ae;
        2452:    rdata = 32'h00b100b0;
        2453:    rdata = 32'h00b300b2;
        2454:    rdata = 32'h00b500b4;
        2455:    rdata = 32'h00b700b6;
        2456:    rdata = 32'h00b900b8;
        2457:    rdata = 32'h00bb00ba;
        2458:    rdata = 32'h00bd00bc;
        2459:    rdata = 32'h00bf00be;
        2460:    rdata = 32'h00c100c0;
        2461:    rdata = 32'h00c300c2;
        2462:    rdata = 32'h00c500c4;
        2463:    rdata = 32'h00c700c6;
        2464:    rdata = 32'h00c900c8;
        2465:    rdata = 32'h00cb00ca;
        2466:    rdata = 32'h00cd00cc;
        2467:    rdata = 32'h00cf00ce;
        2468:    rdata = 32'h00d100d0;
        2469:    rdata = 32'h00d300d2;
        2470:    rdata = 32'h00d500d4;
        2471:    rdata = 32'h00d700d6;
        2472:    rdata = 32'h00d900d8;
        2473:    rdata = 32'h00db00da;
        2474:    rdata = 32'h00dd00dc;
        2475:    rdata = 32'h00df00de;
        2476:    rdata = 32'h00e100e0;
        2477:    rdata = 32'h00e300e2;
        2478:    rdata = 32'h00e500e4;
        2479:    rdata = 32'h00e700e6;
        2480:    rdata = 32'h00e900e8;
        2481:    rdata = 32'h00eb00ea;
        2482:    rdata = 32'h00ed00ec;
        2483:    rdata = 32'h00ef00ee;
        2484:    rdata = 32'h00f100f0;
        2485:    rdata = 32'h00f300f2;
        2486:    rdata = 32'h00f500f4;
        2487:    rdata = 32'h00f700f6;
        2488:    rdata = 32'h00f900f8;
        2489:    rdata = 32'h00fb00fa;
        2490:    rdata = 32'h00fd00fc;
        2491:    rdata = 32'h00ff00fe;
        2492:    rdata = 32'h04010400;
        2493:    rdata = 32'h04030402;
        2494:    rdata = 32'h04050404;
        2495:    rdata = 32'h04070406;
        2496:    rdata = 32'h04090408;
        2497:    rdata = 32'h040b040a;
        2498:    rdata = 32'h040d040c;
        2499:    rdata = 32'h040f040e;
        2500:    rdata = 32'h04110410;
        2501:    rdata = 32'h04130412;
        2502:    rdata = 32'h04150414;
        2503:    rdata = 32'h04170416;
        2504:    rdata = 32'h04190418;
        2505:    rdata = 32'h041b041a;
        2506:    rdata = 32'h041d041c;
        2507:    rdata = 32'h041f041e;
        2508:    rdata = 32'h04210420;
        2509:    rdata = 32'h04230422;
        2510:    rdata = 32'h04250424;
        2511:    rdata = 32'h04270426;
        2512:    rdata = 32'h04290428;
        2513:    rdata = 32'h042b042a;
        2514:    rdata = 32'h042d042c;
        2515:    rdata = 32'h042f042e;
        2516:    rdata = 32'h04310430;
        2517:    rdata = 32'h04330432;
        2518:    rdata = 32'h04350434;
        2519:    rdata = 32'h04370436;
        2520:    rdata = 32'h04390438;
        2521:    rdata = 32'h043b043a;
        2522:    rdata = 32'h043d043c;
        2523:    rdata = 32'h043f043e;
        2524:    rdata = 32'h04410440;
        2525:    rdata = 32'h04430442;
        2526:    rdata = 32'h04450444;
        2527:    rdata = 32'h04470446;
        2528:    rdata = 32'h04490448;
        2529:    rdata = 32'h044b044a;
        2530:    rdata = 32'h044d044c;
        2531:    rdata = 32'h044f044e;
        2532:    rdata = 32'h04510450;
        2533:    rdata = 32'h04530452;
        2534:    rdata = 32'h04550454;
        2535:    rdata = 32'h04570456;
        2536:    rdata = 32'h04590458;
        2537:    rdata = 32'h045b045a;
        2538:    rdata = 32'h045d045c;
        2539:    rdata = 32'h045f045e;
        2540:    rdata = 32'h04610460;
        2541:    rdata = 32'h04630462;
        2542:    rdata = 32'h04650464;
        2543:    rdata = 32'h04670466;
        2544:    rdata = 32'h04690468;
        2545:    rdata = 32'h046b046a;
        2546:    rdata = 32'h046d046c;
        2547:    rdata = 32'h046f046e;
        2548:    rdata = 32'h04710470;
        2549:    rdata = 32'h04730472;
        2550:    rdata = 32'h04750474;
        2551:    rdata = 32'h04770476;
        2552:    rdata = 32'h04790478;
        2553:    rdata = 32'h047b047a;
        2554:    rdata = 32'h047d047c;
        2555:    rdata = 32'h047f047e;
        2556:    rdata = 32'h04810480;
        2557:    rdata = 32'h04830482;
        2558:    rdata = 32'h04850484;
        2559:    rdata = 32'h04870486;
        2560:    rdata = 32'h04890488;
        2561:    rdata = 32'h048b048a;
        2562:    rdata = 32'h048d048c;
        2563:    rdata = 32'h048f048e;
        2564:    rdata = 32'h04910490;
        2565:    rdata = 32'h04930492;
        2566:    rdata = 32'h04950494;
        2567:    rdata = 32'h04970496;
        2568:    rdata = 32'h04990498;
        2569:    rdata = 32'h049b049a;
        2570:    rdata = 32'h049d049c;
        2571:    rdata = 32'h049f049e;
        2572:    rdata = 32'h04a104a0;
        2573:    rdata = 32'h04a304a2;
        2574:    rdata = 32'h04a504a4;
        2575:    rdata = 32'h04a704a6;
        2576:    rdata = 32'h04a904a8;
        2577:    rdata = 32'h04ab04aa;
        2578:    rdata = 32'h04ad04ac;
        2579:    rdata = 32'h04af04ae;
        2580:    rdata = 32'h04b104b0;
        2581:    rdata = 32'h04b304b2;
        2582:    rdata = 32'h04b504b4;
        2583:    rdata = 32'h04b704b6;
        2584:    rdata = 32'h04b904b8;
        2585:    rdata = 32'h04bb04ba;
        2586:    rdata = 32'h04bd04bc;
        2587:    rdata = 32'h04bf04be;
        2588:    rdata = 32'h04c104c0;
        2589:    rdata = 32'h04c304c2;
        2590:    rdata = 32'h04c504c4;
        2591:    rdata = 32'h04c704c6;
        2592:    rdata = 32'h04c904c8;
        2593:    rdata = 32'h04cb04ca;
        2594:    rdata = 32'h04cd04cc;
        2595:    rdata = 32'h04cf04ce;
        2596:    rdata = 32'h04d104d0;
        2597:    rdata = 32'h04d304d2;
        2598:    rdata = 32'h04d504d4;
        2599:    rdata = 32'h04d704d6;
        2600:    rdata = 32'h04d904d8;
        2601:    rdata = 32'h04db04da;
        2602:    rdata = 32'h04dd04dc;
        2603:    rdata = 32'h04df04de;
        2604:    rdata = 32'h04e104e0;
        2605:    rdata = 32'h04e304e2;
        2606:    rdata = 32'h04e504e4;
        2607:    rdata = 32'h04e704e6;
        2608:    rdata = 32'h04e904e8;
        2609:    rdata = 32'h04eb04ea;
        2610:    rdata = 32'h04ed04ec;
        2611:    rdata = 32'h04ef04ee;
        2612:    rdata = 32'h04f104f0;
        2613:    rdata = 32'h04f304f2;
        2614:    rdata = 32'h04f504f4;
        2615:    rdata = 32'h04f704f6;
        2616:    rdata = 32'h04f904f8;
        2617:    rdata = 32'h04fb04fa;
        2618:    rdata = 32'h04fd04fc;
        2619:    rdata = 32'h04ff04fe;
        2620:    rdata = 32'h0002c000;
        2621:    rdata = 32'h0003c000;
        2622:    rdata = 32'hc00002c0;
        2623:    rdata = 32'h02c00003;
        2624:    rdata = 32'h0003c000;
        2625:    rdata = 32'hc00002c0;
        2626:    rdata = 32'h02c00003;
        2627:    rdata = 32'h0003c000;
        2628:    rdata = 32'hc00002c0;
        2629:    rdata = 32'h02c00003;
        2630:    rdata = 32'h0003c000;
        2631:    rdata = 32'hc00002c0;
        2632:    rdata = 32'h02c00003;
        2633:    rdata = 32'h0003c000;
        2634:    rdata = 32'hc00002c0;
        2635:    rdata = 32'h02c00003;
        2636:    rdata = 32'h0003c000;
        2637:    rdata = 32'hc00002c0;
        2638:    rdata = 32'h02c00003;
        2639:    rdata = 32'h0003c000;
        2640:    rdata = 32'hc00002c0;
        2641:    rdata = 32'h02c00003;
        2642:    rdata = 32'h0003c000;
        2643:    rdata = 32'hc00002c0;
        2644:    rdata = 32'h02c00003;
        2645:    rdata = 32'h00042000;
        2646:    rdata = 32'h0002c000;
        2647:    rdata = 32'h0005c000;
        2648:    rdata = 32'hc00004c0;
        2649:    rdata = 32'h04c00005;
        2650:    rdata = 32'h0005c000;
        2651:    rdata = 32'hc00004c0;
        2652:    rdata = 32'h04c00005;
        2653:    rdata = 32'h0005c000;
        2654:    rdata = 32'hc00004c0;
        2655:    rdata = 32'h04c00005;
        2656:    rdata = 32'h0005c000;
        2657:    rdata = 32'hc00004c0;
        2658:    rdata = 32'h04c00005;
        2659:    rdata = 32'h0005c000;
        2660:    rdata = 32'hc00004c0;
        2661:    rdata = 32'h04c00005;
        2662:    rdata = 32'h0005c000;
        2663:    rdata = 32'hc00004c0;
        2664:    rdata = 32'h04c00005;
        2665:    rdata = 32'h0005c000;
        2666:    rdata = 32'hc00004c0;
        2667:    rdata = 32'h04c00005;
        2668:    rdata = 32'h0005c000;
        2669:    rdata = 32'hc00004c0;
        2670:    rdata = 32'h04c00005;
        2671:    rdata = 32'h00042000;
        2672:    rdata = 32'h0003c000;
        2673:    rdata = 32'h200002c0;
        2674:    rdata = 32'h00000000;
        2675:    rdata = 32'h0005c000;
        2676:    rdata = 32'h200004c0;
        2677:    rdata = 32'h00000000;
        2678:    rdata = 32'h0020c000;
        2679:    rdata = 32'h200000c0;
        2680:    rdata = 32'h00000000;
        2681:    rdata = 32'h0008c000;
        2682:    rdata = 32'h200000c0;
        2683:    rdata = 32'h00000000;
        2684:    rdata = 32'h72616568;
        2685:    rdata = 32'h61656274;
        2686:    rdata = 32'h00000a74;
        2687:    rdata = 32'h706c6568;
        2688:    rdata = 32'h20202020;
        2689:    rdata = 32'h20202020;
        2690:    rdata = 32'h20202020;
        2691:    rdata = 32'h20202020;
        2692:    rdata = 32'h20202020;
        2693:    rdata = 32'h20202020;
        2694:    rdata = 32'h20202020;
        2695:    rdata = 32'h202d2020;
        2696:    rdata = 32'h6e697270;
        2697:    rdata = 32'h68742074;
        2698:    rdata = 32'h6d207369;
        2699:    rdata = 32'h61737365;
        2700:    rdata = 32'h720a6567;
        2701:    rdata = 32'h74657365;
        2702:    rdata = 32'h20202020;
        2703:    rdata = 32'h20202020;
        2704:    rdata = 32'h20202020;
        2705:    rdata = 32'h20202020;
        2706:    rdata = 32'h20202020;
        2707:    rdata = 32'h20202020;
        2708:    rdata = 32'h20202020;
        2709:    rdata = 32'h72202d20;
        2710:    rdata = 32'h74657365;
        2711:    rdata = 32'h636f7320;
        2712:    rdata = 32'h6e69700a;
        2713:    rdata = 32'h20202067;
        2714:    rdata = 32'h20202020;
        2715:    rdata = 32'h20202020;
        2716:    rdata = 32'h20202020;
        2717:    rdata = 32'h20202020;
        2718:    rdata = 32'h20202020;
        2719:    rdata = 32'h20202020;
        2720:    rdata = 32'h2d202020;
        2721:    rdata = 32'h6e657320;
        2722:    rdata = 32'h70222064;
        2723:    rdata = 32'h22676e69;
        2724:    rdata = 32'h206f7420;
        2725:    rdata = 32'h20656874;
        2726:    rdata = 32'h74736f68;
        2727:    rdata = 32'h7465730a;
        2728:    rdata = 32'h6970675f;
        2729:    rdata = 32'h69645f6f;
        2730:    rdata = 32'h74636572;
        2731:    rdata = 32'h206e6f69;
        2732:    rdata = 32'h6e69703c;
        2733:    rdata = 32'h695b203e;
        2734:    rdata = 32'h756f7c6e;
        2735:    rdata = 32'h2d205d74;
        2736:    rdata = 32'h74657320;
        2737:    rdata = 32'h69706720;
        2738:    rdata = 32'h6970206f;
        2739:    rdata = 32'h6964206e;
        2740:    rdata = 32'h74636572;
        2741:    rdata = 32'h0a6e6f69;
        2742:    rdata = 32'h5f746567;
        2743:    rdata = 32'h6f697067;
        2744:    rdata = 32'h7269645f;
        2745:    rdata = 32'h69746365;
        2746:    rdata = 32'h3c206e6f;
        2747:    rdata = 32'h3e6e6970;
        2748:    rdata = 32'h20202020;
        2749:    rdata = 32'h20202020;
        2750:    rdata = 32'h202d2020;
        2751:    rdata = 32'h20746567;
        2752:    rdata = 32'h6f697067;
        2753:    rdata = 32'h6e697020;
        2754:    rdata = 32'h72696420;
        2755:    rdata = 32'h69746365;
        2756:    rdata = 32'h730a6e6f;
        2757:    rdata = 32'h675f7465;
        2758:    rdata = 32'h206f6970;
        2759:    rdata = 32'h6e69703c;
        2760:    rdata = 32'h763c203e;
        2761:    rdata = 32'h65756c61;
        2762:    rdata = 32'h2020203e;
        2763:    rdata = 32'h20202020;
        2764:    rdata = 32'h20202020;
        2765:    rdata = 32'h73202d20;
        2766:    rdata = 32'h67207465;
        2767:    rdata = 32'h206f6970;
        2768:    rdata = 32'h0a6e6970;
        2769:    rdata = 32'h5f746567;
        2770:    rdata = 32'h6f697067;
        2771:    rdata = 32'h69703c20;
        2772:    rdata = 32'h20203e6e;
        2773:    rdata = 32'h20202020;
        2774:    rdata = 32'h20202020;
        2775:    rdata = 32'h20202020;
        2776:    rdata = 32'h20202020;
        2777:    rdata = 32'h202d2020;
        2778:    rdata = 32'h20746567;
        2779:    rdata = 32'h6f697067;
        2780:    rdata = 32'h6e697020;
        2781:    rdata = 32'h7465730a;
        2782:    rdata = 32'h6165685f;
        2783:    rdata = 32'h65627472;
        2784:    rdata = 32'h3c207461;
        2785:    rdata = 32'h69726570;
        2786:    rdata = 32'h5b20646f;
        2787:    rdata = 32'h3e5d736d;
        2788:    rdata = 32'h20202020;
        2789:    rdata = 32'h2d202020;
        2790:    rdata = 32'h74657320;
        2791:    rdata = 32'h61656820;
        2792:    rdata = 32'h65627472;
        2793:    rdata = 32'h630a7461;
        2794:    rdata = 32'h75636c61;
        2795:    rdata = 32'h6574616c;
        2796:    rdata = 32'h72613c20;
        2797:    rdata = 32'h203e3167;
        2798:    rdata = 32'h2d7c2b5b;
        2799:    rdata = 32'h2f7c2a7c;
        2800:    rdata = 32'h613c205d;
        2801:    rdata = 32'h3e326772;
        2802:    rdata = 32'h70202d20;
        2803:    rdata = 32'h6f667265;
        2804:    rdata = 32'h63206d72;
        2805:    rdata = 32'h75636c61;
        2806:    rdata = 32'h6974616c;
        2807:    rdata = 32'h730a6e6f;
        2808:    rdata = 32'h705f7465;
        2809:    rdata = 32'h6f635f6d;
        2810:    rdata = 32'h6f72746e;
        2811:    rdata = 32'h72656c6c;
        2812:    rdata = 32'h646f6d5f;
        2813:    rdata = 32'h6d3c2065;
        2814:    rdata = 32'h3e65646f;
        2815:    rdata = 32'h20202020;
        2816:    rdata = 32'h73202d20;
        2817:    rdata = 32'h70207465;
        2818:    rdata = 32'h6f63206d;
        2819:    rdata = 32'h6f72746e;
        2820:    rdata = 32'h72656c6c;
        2821:    rdata = 32'h646f6d20;
        2822:    rdata = 32'h2d200a65;
        2823:    rdata = 32'h63636120;
        2824:    rdata = 32'h72656c65;
        2825:    rdata = 32'h64657461;
        2826:    rdata = 32'h202d200a;
        2827:    rdata = 32'h72706f63;
        2828:    rdata = 32'h7365636f;
        2829:    rdata = 32'h0a646573;
        2830:    rdata = 32'h64202d20;
        2831:    rdata = 32'h63657269;
        2832:    rdata = 32'h65720a74;
        2833:    rdata = 32'h6d5f6461;
        2834:    rdata = 32'h69727461;
        2835:    rdata = 32'h20202078;
        2836:    rdata = 32'h20202020;
        2837:    rdata = 32'h20202020;
        2838:    rdata = 32'h20202020;
        2839:    rdata = 32'h20202020;
        2840:    rdata = 32'h20202020;
        2841:    rdata = 32'h6572202d;
        2842:    rdata = 32'h6d206461;
        2843:    rdata = 32'h69727461;
        2844:    rdata = 32'h61630a78;
        2845:    rdata = 32'h7262696c;
        2846:    rdata = 32'h5f657461;
        2847:    rdata = 32'h7274616d;
        2848:    rdata = 32'h20207869;
        2849:    rdata = 32'h20202020;
        2850:    rdata = 32'h20202020;
        2851:    rdata = 32'h20202020;
        2852:    rdata = 32'h20202020;
        2853:    rdata = 32'h6163202d;
        2854:    rdata = 32'h7262696c;
        2855:    rdata = 32'h20657461;
        2856:    rdata = 32'h65786970;
        2857:    rdata = 32'h6f20736c;
        2858:    rdata = 32'h65736666;
        2859:    rdata = 32'h740a7374;
        2860:    rdata = 32'h5f747365;
        2861:    rdata = 32'h7274616d;
        2862:    rdata = 32'h775f7869;
        2863:    rdata = 32'h65746972;
        2864:    rdata = 32'h6165725f;
        2865:    rdata = 32'h20202064;
        2866:    rdata = 32'h20202020;
        2867:    rdata = 32'h20202020;
        2868:    rdata = 32'h65202d20;
        2869:    rdata = 32'h75636578;
        2870:    rdata = 32'h6d206574;
        2871:    rdata = 32'h69727461;
        2872:    rdata = 32'h72772078;
        2873:    rdata = 32'h5f657469;
        2874:    rdata = 32'h64616572;
        2875:    rdata = 32'h73657420;
        2876:    rdata = 32'h00000a74;
        2877:    rdata = 32'h6f727265;
        2878:    rdata = 32'h6f203a72;
        2879:    rdata = 32'h61726570;
        2880:    rdata = 32'h6e6f6974;
        2881:    rdata = 32'h746f6e20;
        2882:    rdata = 32'h70757320;
        2883:    rdata = 32'h74726f70;
        2884:    rdata = 32'h000a6465;
        2885:    rdata = 32'h676e6970;
        2886:    rdata = 32'h0000000a;
        2887:    rdata = 32'h6f727265;
        2888:    rdata = 32'h6d203a72;
        2889:    rdata = 32'h69737369;
        2890:    rdata = 32'h6120676e;
        2891:    rdata = 32'h6d756772;
        2892:    rdata = 32'h28746e65;
        2893:    rdata = 32'h000a2973;
        2894:    rdata = 32'h6f727265;
        2895:    rdata = 32'h69203a72;
        2896:    rdata = 32'h6c61766e;
        2897:    rdata = 32'h61206469;
        2898:    rdata = 32'h6d756772;
        2899:    rdata = 32'h28746e65;
        2900:    rdata = 32'h74202973;
        2901:    rdata = 32'h28657079;
        2902:    rdata = 32'h000a2973;
        2903:    rdata = 32'h00006e69;
        2904:    rdata = 32'h0074756f;
        2905:    rdata = 32'h6f727265;
        2906:    rdata = 32'h69203a72;
        2907:    rdata = 32'h6c61766e;
        2908:    rdata = 32'h64206469;
        2909:    rdata = 32'h63657269;
        2910:    rdata = 32'h6e6f6974;
        2911:    rdata = 32'h0000000a;
        2912:    rdata = 32'h6f727265;
        2913:    rdata = 32'h6d203a72;
        2914:    rdata = 32'h69737369;
        2915:    rdata = 32'h6120676e;
        2916:    rdata = 32'h6d756772;
        2917:    rdata = 32'h0a746e65;
        2918:    rdata = 32'h00000000;
        2919:    rdata = 32'h6f727265;
        2920:    rdata = 32'h69203a72;
        2921:    rdata = 32'h6c61766e;
        2922:    rdata = 32'h61206469;
        2923:    rdata = 32'h6d756772;
        2924:    rdata = 32'h20746e65;
        2925:    rdata = 32'h65707974;
        2926:    rdata = 32'h0000000a;
        2927:    rdata = 32'h6f727265;
        2928:    rdata = 32'h64203a72;
        2929:    rdata = 32'h73697669;
        2930:    rdata = 32'h206e6f69;
        2931:    rdata = 32'h7a207962;
        2932:    rdata = 32'h0a6f7265;
        2933:    rdata = 32'h00000000;
        2934:    rdata = 32'h6f727265;
        2935:    rdata = 32'h75203a72;
        2936:    rdata = 32'h6365726e;
        2937:    rdata = 32'h696e676f;
        2938:    rdata = 32'h2064657a;
        2939:    rdata = 32'h7265706f;
        2940:    rdata = 32'h6f697461;
        2941:    rdata = 32'h00000a6e;
        2942:    rdata = 32'h65636361;
        2943:    rdata = 32'h6172656c;
        2944:    rdata = 32'h00646574;
        2945:    rdata = 32'h72706f63;
        2946:    rdata = 32'h7365636f;
        2947:    rdata = 32'h00646573;
        2948:    rdata = 32'h65726964;
        2949:    rdata = 32'h00007463;
        2950:    rdata = 32'h6f727265;
        2951:    rdata = 32'h69203a72;
        2952:    rdata = 32'h6c61766e;
        2953:    rdata = 32'h63206469;
        2954:    rdata = 32'h72746e6f;
        2955:    rdata = 32'h656c6c6f;
        2956:    rdata = 32'h6f6d2072;
        2957:    rdata = 32'h000a6564;
        2958:    rdata = 32'h746e6f63;
        2959:    rdata = 32'h6c6c6f72;
        2960:    rdata = 32'h6d207265;
        2961:    rdata = 32'h2065646f;
        2962:    rdata = 32'h61647075;
        2963:    rdata = 32'h0a646574;
        2964:    rdata = 32'h00000000;
        2965:    rdata = 32'h64616572;
        2966:    rdata = 32'h5f74756f;
        2967:    rdata = 32'h656d6974;
        2968:    rdata = 32'h00000000;
        2969:    rdata = 32'h7366666f;
        2970:    rdata = 32'h63207465;
        2971:    rdata = 32'h62696c61;
        2972:    rdata = 32'h69746172;
        2973:    rdata = 32'h64206e6f;
        2974:    rdata = 32'h0a656e6f;
        2975:    rdata = 32'h00000000;
        2976:    rdata = 32'h696c6163;
        2977:    rdata = 32'h74617262;
        2978:    rdata = 32'h5f6e6f69;
        2979:    rdata = 32'h656d6974;
        2980:    rdata = 32'h00000000;
        2981:    rdata = 32'h73736170;
        2982:    rdata = 32'h00006465;
        2983:    rdata = 32'h6c696166;
        2984:    rdata = 32'h00006465;
        2985:    rdata = 32'h74736574;
        2986:    rdata = 32'h00000020;
        2987:    rdata = 32'h0000203e;
        2988:    rdata = 32'h6f727265;
        2989:    rdata = 32'h75203a72;
        2990:    rdata = 32'h6365726e;
        2991:    rdata = 32'h696e676f;
        2992:    rdata = 32'h2064657a;
        2993:    rdata = 32'h6d6d6f63;
        2994:    rdata = 32'h3a646e61;
        2995:    rdata = 32'h00002220;
        2996:    rdata = 32'h65202e22;
        2997:    rdata = 32'h75636578;
        2998:    rdata = 32'h22206574;
        2999:    rdata = 32'h706c6568;
        3000:    rdata = 32'h6f742022;
        3001:    rdata = 32'h74656720;
        3002:    rdata = 32'h70757320;
        3003:    rdata = 32'h74726f70;
        3004:    rdata = 32'h63206465;
        3005:    rdata = 32'h616d6d6f;
        3006:    rdata = 32'h2073646e;
        3007:    rdata = 32'h7473696c;
        3008:    rdata = 32'h0000000a;
        3009:    rdata = 32'h6f727265;
        3010:    rdata = 32'h63203a72;
        3011:    rdata = 32'h616d6d6f;
        3012:    rdata = 32'h6620646e;
        3013:    rdata = 32'h656c6961;
        3014:    rdata = 32'h00000a64;
        3015:    rdata = 32'h706c6568;
        3016:    rdata = 32'h00000000;
        3017:    rdata = 32'h65736572;
        3018:    rdata = 32'h00000074;
        3019:    rdata = 32'h676e6970;
        3020:    rdata = 32'h00000000;
        3021:    rdata = 32'h5f746573;
        3022:    rdata = 32'h6f697067;
        3023:    rdata = 32'h7269645f;
        3024:    rdata = 32'h69746365;
        3025:    rdata = 32'h00006e6f;
        3026:    rdata = 32'h5f746567;
        3027:    rdata = 32'h6f697067;
        3028:    rdata = 32'h7269645f;
        3029:    rdata = 32'h69746365;
        3030:    rdata = 32'h00006e6f;
        3031:    rdata = 32'h5f746573;
        3032:    rdata = 32'h6f697067;
        3033:    rdata = 32'h00000000;
        3034:    rdata = 32'h5f746567;
        3035:    rdata = 32'h6f697067;
        3036:    rdata = 32'h00000000;
        3037:    rdata = 32'h5f746573;
        3038:    rdata = 32'h72616568;
        3039:    rdata = 32'h61656274;
        3040:    rdata = 32'h00000074;
        3041:    rdata = 32'h636c6163;
        3042:    rdata = 32'h74616c75;
        3043:    rdata = 32'h00000065;
        3044:    rdata = 32'h5f746573;
        3045:    rdata = 32'h635f6d70;
        3046:    rdata = 32'h72746e6f;
        3047:    rdata = 32'h656c6c6f;
        3048:    rdata = 32'h6f6d5f72;
        3049:    rdata = 32'h00006564;
        3050:    rdata = 32'h64616572;
        3051:    rdata = 32'h74616d5f;
        3052:    rdata = 32'h00786972;
        3053:    rdata = 32'h696c6163;
        3054:    rdata = 32'h74617262;
        3055:    rdata = 32'h616d5f65;
        3056:    rdata = 32'h78697274;
        3057:    rdata = 32'h00000000;
        3058:    rdata = 32'h74736574;
        3059:    rdata = 32'h74616d5f;
        3060:    rdata = 32'h5f786972;
        3061:    rdata = 32'h74697277;
        3062:    rdata = 32'h65725f65;
        3063:    rdata = 32'h00006461;
        3064:    rdata = 32'h6d6d6f63;
        3065:    rdata = 32'h5f646e61;
        3066:    rdata = 32'h65746e69;
        3067:    rdata = 32'h65727072;
        3068:    rdata = 32'h20726574;
        3069:    rdata = 32'h72617473;
        3070:    rdata = 32'h0a646574;
        3071:    rdata = 32'h00000000;
        3072:    rdata = 32'h0000203a;
        3073:    rdata = 32'h00002820;
        3074:    rdata = 32'h00203a29;
        3075:    rdata = 32'h6f636e69;
        3076:    rdata = 32'h63657272;
        3077:    rdata = 32'h61762074;
        3078:    rdata = 32'h2e65756c;
        3079:    rdata = 32'h79727420;
        3080:    rdata = 32'h61676120;
        3081:    rdata = 32'h000a6e69;
        default: rdata = 32'h00000000;
    endcase
end
endmodule
