/**
 * Copyright (C) 2020  AGH University of Science and Technology
 *
 * This program is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with this program.  If not, see <https://www.gnu.org/licenses/>.
 */

module boot_mem (
    output logic [31:0] rdata,
    input logic [31:0] addr
);

/**
 * Module internal logic
 */

always_comb begin
    case (addr[13:2])
           0:    rdata = 32'h08c0006f;
           1:    rdata = 32'h0880006f;
           2:    rdata = 32'h0840006f;
           3:    rdata = 32'h0800006f;
           4:    rdata = 32'h07c0006f;
           5:    rdata = 32'h0780006f;
           6:    rdata = 32'h0740006f;
           7:    rdata = 32'h0700006f;
           8:    rdata = 32'h06c0006f;
           9:    rdata = 32'h0680006f;
          10:    rdata = 32'h0640006f;
          11:    rdata = 32'h0600006f;
          12:    rdata = 32'h05c0006f;
          13:    rdata = 32'h0580006f;
          14:    rdata = 32'h0540006f;
          15:    rdata = 32'h0500006f;
          16:    rdata = 32'h04c0006f;
          17:    rdata = 32'h0480006f;
          18:    rdata = 32'h0440006f;
          19:    rdata = 32'h0400006f;
          20:    rdata = 32'h03c0006f;
          21:    rdata = 32'h0380006f;
          22:    rdata = 32'h0340006f;
          23:    rdata = 32'h0300006f;
          24:    rdata = 32'h02c0006f;
          25:    rdata = 32'h0280006f;
          26:    rdata = 32'h0240006f;
          27:    rdata = 32'h0200006f;
          28:    rdata = 32'h01c0006f;
          29:    rdata = 32'h0180006f;
          30:    rdata = 32'h0140006f;
          31:    rdata = 32'h0100006f;
          32:    rdata = 32'h0100006f;
          33:    rdata = 32'h0080006f;
          34:    rdata = 32'h0040006f;
          35:    rdata = 32'h0000006f;
          36:    rdata = 32'h00000093;
          37:    rdata = 32'h00000113;
          38:    rdata = 32'h00000193;
          39:    rdata = 32'h00000213;
          40:    rdata = 32'h00000293;
          41:    rdata = 32'h00000313;
          42:    rdata = 32'h00000393;
          43:    rdata = 32'h00000413;
          44:    rdata = 32'h00000493;
          45:    rdata = 32'h00000513;
          46:    rdata = 32'h00000593;
          47:    rdata = 32'h00000613;
          48:    rdata = 32'h00000693;
          49:    rdata = 32'h00000713;
          50:    rdata = 32'h00000793;
          51:    rdata = 32'h00000813;
          52:    rdata = 32'h00000893;
          53:    rdata = 32'h00000913;
          54:    rdata = 32'h00000993;
          55:    rdata = 32'h00000a13;
          56:    rdata = 32'h00000a93;
          57:    rdata = 32'h00000b13;
          58:    rdata = 32'h00000b93;
          59:    rdata = 32'h00000c13;
          60:    rdata = 32'h00000c93;
          61:    rdata = 32'h00000d13;
          62:    rdata = 32'h00000d93;
          63:    rdata = 32'h00000e13;
          64:    rdata = 32'h00000e93;
          65:    rdata = 32'h00000f13;
          66:    rdata = 32'h00000f93;
          67:    rdata = 32'h00104117;
          68:    rdata = 32'hef410113;
          69:    rdata = 32'h00100297;
          70:    rdata = 32'heec28293;
          71:    rdata = 32'h00100317;
          72:    rdata = 32'hf0c30313;
          73:    rdata = 32'h0062d863;
          74:    rdata = 32'h0002a023;
          75:    rdata = 32'h00428293;
          76:    rdata = 32'hfe535ce3;
          77:    rdata = 32'h00001297;
          78:    rdata = 32'h0fc28293;
          79:    rdata = 32'h00100317;
          80:    rdata = 32'hec430313;
          81:    rdata = 32'h00100397;
          82:    rdata = 32'hebc38393;
          83:    rdata = 32'h00735c63;
          84:    rdata = 32'h0002ae03;
          85:    rdata = 32'h01c32023;
          86:    rdata = 32'h00428293;
          87:    rdata = 32'h00430313;
          88:    rdata = 32'hfe7348e3;
          89:    rdata = 32'h00001297;
          90:    rdata = 32'hfc428293;
          91:    rdata = 32'h00001317;
          92:    rdata = 32'hfcc30313;
          93:    rdata = 32'h0062da63;
          94:    rdata = 32'h0002a783;
          95:    rdata = 32'h000780e7;
          96:    rdata = 32'h00428293;
          97:    rdata = 32'hfe62cae3;
          98:    rdata = 32'h00000513;
          99:    rdata = 32'h00000593;
         100:    rdata = 32'h621000ef;
         101:    rdata = 32'h65c16611;
         102:    rdata = 32'h7179a585;
         103:    rdata = 32'h4581d226;
         104:    rdata = 32'h051784aa;
         105:    rdata = 32'h05130010;
         106:    rdata = 32'hd606e7e5;
         107:    rdata = 32'hce4ed422;
         108:    rdata = 32'hd04acc52;
         109:    rdata = 32'h23b000ef;
         110:    rdata = 32'h05174585;
         111:    rdata = 32'h05130010;
         112:    rdata = 32'h00efe665;
         113:    rdata = 32'h458d2390;
         114:    rdata = 32'h00100517;
         115:    rdata = 32'he5850513;
         116:    rdata = 32'h243000ef;
         117:    rdata = 32'h09974401;
         118:    rdata = 32'h89930010;
         119:    rdata = 32'h4a11e4a9;
         120:    rdata = 32'h2d158526;
         121:    rdata = 32'h02a47363;
         122:    rdata = 32'h854e4901;
         123:    rdata = 32'h2c1000ef;
         124:    rdata = 32'h97ca007c;
         125:    rdata = 32'h00a78023;
         126:    rdata = 32'h18e30905;
         127:    rdata = 32'h4632ff49;
         128:    rdata = 32'h852685a2;
         129:    rdata = 32'h04112519;
         130:    rdata = 32'h50b2bfe1;
         131:    rdata = 32'h54925422;
         132:    rdata = 32'h49f25902;
         133:    rdata = 32'h61454a62;
         134:    rdata = 32'h71398082;
         135:    rdata = 32'hd452d84a;
         136:    rdata = 32'h3b9ad937;
         137:    rdata = 32'h05178a2a;
         138:    rdata = 32'h05130010;
         139:    rdata = 32'hdc22dda5;
         140:    rdata = 32'hd64eda26;
         141:    rdata = 32'hce5ed256;
         142:    rdata = 32'hd05ade06;
         143:    rdata = 32'h0913cc62;
         144:    rdata = 32'h2be1a009;
         145:    rdata = 32'h3433992a;
         146:    rdata = 32'h942e00a9;
         147:    rdata = 32'h44814981;
         148:    rdata = 32'h00100a97;
         149:    rdata = 32'hdd4a8a93;
         150:    rdata = 32'h00100b97;
         151:    rdata = 32'hda8b8b93;
         152:    rdata = 32'h2b558552;
         153:    rdata = 32'h04a9f563;
         154:    rdata = 32'h00c10b13;
         155:    rdata = 32'h00448c13;
         156:    rdata = 32'h00ef8556;
         157:    rdata = 32'he90935b0;
         158:    rdata = 32'h2345855e;
         159:    rdata = 32'hfe85eae3;
         160:    rdata = 32'h00b41463;
         161:    rdata = 32'hff2566e3;
         162:    rdata = 32'h00ef8556;
         163:    rdata = 32'hc10d3430;
         164:    rdata = 32'h00ef8556;
         165:    rdata = 32'h00233530;
         166:    rdata = 32'h048500ab;
         167:    rdata = 32'h99e30b05;
         168:    rdata = 32'h4632fd84;
         169:    rdata = 32'h855285ce;
         170:    rdata = 32'h0991238d;
         171:    rdata = 32'h4481bf55;
         172:    rdata = 32'h546250f2;
         173:    rdata = 32'h59b25942;
         174:    rdata = 32'h5a925a22;
         175:    rdata = 32'h4bf25b02;
         176:    rdata = 32'h85264c62;
         177:    rdata = 32'h612154d2;
         178:    rdata = 32'h00238082;
         179:    rdata = 32'h460100b5;
         180:    rdata = 32'h00100517;
         181:    rdata = 32'hd4850513;
         182:    rdata = 32'h7880006f;
         183:    rdata = 32'hc4221141;
         184:    rdata = 32'h0513842a;
         185:    rdata = 32'hc6060fa0;
         186:    rdata = 32'h45832a01;
         187:    rdata = 32'h46050004;
         188:    rdata = 32'h00100517;
         189:    rdata = 32'hd2850513;
         190:    rdata = 32'h790000ef;
         191:    rdata = 32'h0fa00513;
         192:    rdata = 32'h458328e5;
         193:    rdata = 32'h05170004;
         194:    rdata = 32'h05130010;
         195:    rdata = 32'h4601d125;
         196:    rdata = 32'h778000ef;
         197:    rdata = 32'h40b24422;
         198:    rdata = 32'h0fa00513;
         199:    rdata = 32'ha8e90141;
         200:    rdata = 32'hc4221141;
         201:    rdata = 32'h0513842a;
         202:    rdata = 32'hc6060fa0;
         203:    rdata = 32'h458320f1;
         204:    rdata = 32'h46050004;
         205:    rdata = 32'h00100517;
         206:    rdata = 32'hce450513;
         207:    rdata = 32'h74c000ef;
         208:    rdata = 32'h0fa00513;
         209:    rdata = 32'h45832855;
         210:    rdata = 32'h46010004;
         211:    rdata = 32'h00100517;
         212:    rdata = 32'hccc50513;
         213:    rdata = 32'h734000ef;
         214:    rdata = 32'h0fa00513;
         215:    rdata = 32'h45832871;
         216:    rdata = 32'h46050004;
         217:    rdata = 32'h00100517;
         218:    rdata = 32'hcb450513;
         219:    rdata = 32'h71c000ef;
         220:    rdata = 32'h0fa00513;
         221:    rdata = 32'h45832051;
         222:    rdata = 32'h46010004;
         223:    rdata = 32'h00100517;
         224:    rdata = 32'hc9c50513;
         225:    rdata = 32'h704000ef;
         226:    rdata = 32'h0fa00513;
         227:    rdata = 32'h442220b5;
         228:    rdata = 32'h051340b2;
         229:    rdata = 32'h01410fa0;
         230:    rdata = 32'h1141a085;
         231:    rdata = 32'h842ac422;
         232:    rdata = 32'h0fa00513;
         233:    rdata = 32'hc606c226;
         234:    rdata = 32'h00100497;
         235:    rdata = 32'hc7048493;
         236:    rdata = 32'h458320a1;
         237:    rdata = 32'h46050004;
         238:    rdata = 32'h25f98526;
         239:    rdata = 32'h0fa00513;
         240:    rdata = 32'h45832825;
         241:    rdata = 32'h85260004;
         242:    rdata = 32'h2d7d4601;
         243:    rdata = 32'h0fa00513;
         244:    rdata = 32'hb7c52025;
         245:    rdata = 32'hc4221141;
         246:    rdata = 32'h0513842a;
         247:    rdata = 32'hc6060fa0;
         248:    rdata = 32'h45832821;
         249:    rdata = 32'h44220004;
         250:    rdata = 32'h460540b2;
         251:    rdata = 32'h00100517;
         252:    rdata = 32'hc2c50513;
         253:    rdata = 32'had490141;
         254:    rdata = 32'h87936785;
         255:    rdata = 32'h05b33887;
         256:    rdata = 32'h051702f5;
         257:    rdata = 32'h05130010;
         258:    rdata = 32'ha929bfe5;
         259:    rdata = 32'h05b34595;
         260:    rdata = 32'h051702b5;
         261:    rdata = 32'h05130010;
         262:    rdata = 32'ha129bee5;
         263:    rdata = 32'hc4221141;
         264:    rdata = 32'h06400613;
         265:    rdata = 32'h0517842a;
         266:    rdata = 32'h05130010;
         267:    rdata = 32'hc606bfe5;
         268:    rdata = 32'h1e7000ef;
         269:    rdata = 32'h852240b2;
         270:    rdata = 32'h01414422;
         271:    rdata = 32'h11418082;
         272:    rdata = 32'h842ac422;
         273:    rdata = 32'h00100517;
         274:    rdata = 32'hbe050513;
         275:    rdata = 32'h00efc606;
         276:    rdata = 32'h40b226b0;
         277:    rdata = 32'h44228522;
         278:    rdata = 32'h80820141;
         279:    rdata = 32'hc4221141;
         280:    rdata = 32'h0517842a;
         281:    rdata = 32'h05130010;
         282:    rdata = 32'hc606bc25;
         283:    rdata = 32'h24d000ef;
         284:    rdata = 32'h852240b2;
         285:    rdata = 32'h01414422;
         286:    rdata = 32'h418c8082;
         287:    rdata = 32'hcc221101;
         288:    rdata = 32'h0048842a;
         289:    rdata = 32'h2c35ce06;
         290:    rdata = 32'h0517004c;
         291:    rdata = 32'h05130010;
         292:    rdata = 32'h00efb9a5;
         293:    rdata = 32'h40f22270;
         294:    rdata = 32'h44628522;
         295:    rdata = 32'h80826105;
         296:    rdata = 32'hc4221141;
         297:    rdata = 32'h0417c606;
         298:    rdata = 32'h04130010;
         299:    rdata = 32'h8522b7e4;
         300:    rdata = 32'h1c7000ef;
         301:    rdata = 32'h40b2fd6d;
         302:    rdata = 32'h01414422;
         303:    rdata = 32'h71758082;
         304:    rdata = 32'hc326c522;
         305:    rdata = 32'hdecec14a;
         306:    rdata = 32'hc706dcd2;
         307:    rdata = 32'h892e84aa;
         308:    rdata = 32'h00100417;
         309:    rdata = 32'hb5440413;
         310:    rdata = 32'h00001a17;
         311:    rdata = 32'hce4a0a13;
         312:    rdata = 32'h00001997;
         313:    rdata = 32'hd3498993;
         314:    rdata = 32'h852285ca;
         315:    rdata = 32'h1cd000ef;
         316:    rdata = 32'h852285d2;
         317:    rdata = 32'h1c5000ef;
         318:    rdata = 32'h8526006c;
         319:    rdata = 32'h00683705;
         320:    rdata = 32'he5112411;
         321:    rdata = 32'h852285ce;
         322:    rdata = 32'h1b1000ef;
         323:    rdata = 32'h0068bff1;
         324:    rdata = 32'h40ba242d;
         325:    rdata = 32'h449a442a;
         326:    rdata = 32'h59f6490a;
         327:    rdata = 32'h61495a66;
         328:    rdata = 32'h07138082;
         329:    rdata = 32'h47830300;
         330:    rdata = 32'h94630005;
         331:    rdata = 32'h050500e7;
         332:    rdata = 32'he391bfdd;
         333:    rdata = 32'h8082157d;
         334:    rdata = 32'h00054703;
         335:    rdata = 32'h02d00793;
         336:    rdata = 32'h00f71363;
         337:    rdata = 32'h47250505;
         338:    rdata = 32'h00054783;
         339:    rdata = 32'hfd078793;
         340:    rdata = 32'h0ff7f793;
         341:    rdata = 32'h00f76863;
         342:    rdata = 32'h00154783;
         343:    rdata = 32'hf7ed0505;
         344:    rdata = 32'h80824505;
         345:    rdata = 32'h80824501;
         346:    rdata = 32'h46a50509;
         347:    rdata = 32'h47834615;
         348:    rdata = 32'h87130005;
         349:    rdata = 32'h7713fd07;
         350:    rdata = 32'hfa630ff7;
         351:    rdata = 32'hf79300e6;
         352:    rdata = 32'h8793fdf7;
         353:    rdata = 32'hf793fbf7;
         354:    rdata = 32'h68630ff7;
         355:    rdata = 32'h478300f6;
         356:    rdata = 32'h05050015;
         357:    rdata = 32'h4505ffe9;
         358:    rdata = 32'h45018082;
         359:    rdata = 32'h87aa8082;
         360:    rdata = 32'h0005c703;
         361:    rdata = 32'h07850585;
         362:    rdata = 32'hfee78fa3;
         363:    rdata = 32'h8082fb75;
         364:    rdata = 32'hc68387aa;
         365:    rdata = 32'h873e0007;
         366:    rdata = 32'hfee50785;
         367:    rdata = 32'h0005c783;
         368:    rdata = 32'h07050585;
         369:    rdata = 32'hfef70fa3;
         370:    rdata = 32'h8082fbf5;
         371:    rdata = 32'h00054783;
         372:    rdata = 32'h0005c703;
         373:    rdata = 32'h00e78763;
         374:    rdata = 32'he963557d;
         375:    rdata = 32'h450500e7;
         376:    rdata = 32'hc7818082;
         377:    rdata = 32'h05850505;
         378:    rdata = 32'h4501b7d5;
         379:    rdata = 32'h87aa8082;
         380:    rdata = 32'h87334501;
         381:    rdata = 32'h470300a7;
         382:    rdata = 32'hc3190007;
         383:    rdata = 32'hbfd50505;
         384:    rdata = 32'h47898082;
         385:    rdata = 32'h02f60c63;
         386:    rdata = 32'h0d634791;
         387:    rdata = 32'h470502f6;
         388:    rdata = 32'h14634781;
         389:    rdata = 32'h079300e6;
         390:    rdata = 32'h46290640;
         391:    rdata = 32'hd733cb8d;
         392:    rdata = 32'h050502f5;
         393:    rdata = 32'h0ff77693;
         394:    rdata = 32'h02f686b3;
         395:    rdata = 32'h03070713;
         396:    rdata = 32'hfee50fa3;
         397:    rdata = 32'h02c7d7b3;
         398:    rdata = 32'hb7cd8d95;
         399:    rdata = 32'h87936789;
         400:    rdata = 32'hbfe17107;
         401:    rdata = 32'h3b9ad7b7;
         402:    rdata = 32'ha0078793;
         403:    rdata = 32'h0023b7f9;
         404:    rdata = 32'h80820005;
         405:    rdata = 32'hb7754605;
         406:    rdata = 32'hcc221101;
         407:    rdata = 32'h842a4611;
         408:    rdata = 32'hce060048;
         409:    rdata = 32'h00483f79;
         410:    rdata = 32'h85aa3d6d;
         411:    rdata = 32'h3f058522;
         412:    rdata = 32'h446240f2;
         413:    rdata = 32'h80826105;
         414:    rdata = 32'h03000793;
         415:    rdata = 32'h76130606;
         416:    rdata = 32'h00230ff6;
         417:    rdata = 32'h079300f5;
         418:    rdata = 32'h00a30780;
         419:    rdata = 32'h482500f5;
         420:    rdata = 32'hc38587b2;
         421:    rdata = 32'h00f5f713;
         422:    rdata = 32'h05770693;
         423:    rdata = 32'h00e86463;
         424:    rdata = 32'h03070693;
         425:    rdata = 32'h00f50733;
         426:    rdata = 32'h00d700a3;
         427:    rdata = 32'h17fd8191;
         428:    rdata = 32'h9532b7cd;
         429:    rdata = 32'h00050123;
         430:    rdata = 32'h46058082;
         431:    rdata = 32'h4611bf75;
         432:    rdata = 32'h1101bf65;
         433:    rdata = 32'hce06cc22;
         434:    rdata = 32'hd563842a;
         435:    rdata = 32'h07130205;
         436:    rdata = 32'h002302d0;
         437:    rdata = 32'h05b300e5;
         438:    rdata = 32'h461140b0;
         439:    rdata = 32'h37150048;
         440:    rdata = 32'h35810048;
         441:    rdata = 32'h051385aa;
         442:    rdata = 32'h3d550014;
         443:    rdata = 32'h446240f2;
         444:    rdata = 32'h80826105;
         445:    rdata = 32'h00484611;
         446:    rdata = 32'h00483729;
         447:    rdata = 32'h85aa351d;
         448:    rdata = 32'hb7e58522;
         449:    rdata = 32'hc4221141;
         450:    rdata = 32'h842ac606;
         451:    rdata = 32'he1153535;
         452:    rdata = 32'h00044703;
         453:    rdata = 32'h03000793;
         454:    rdata = 32'h00f71d63;
         455:    rdata = 32'h00144703;
         456:    rdata = 32'h07800793;
         457:    rdata = 32'h00f71763;
         458:    rdata = 32'h44228522;
         459:    rdata = 32'h014140b2;
         460:    rdata = 32'h40b2bd25;
         461:    rdata = 32'h01414422;
         462:    rdata = 32'h11418082;
         463:    rdata = 32'hc606c422;
         464:    rdata = 32'h3bdd842a;
         465:    rdata = 32'h00044783;
         466:    rdata = 32'h0693c91d;
         467:    rdata = 32'h470102d0;
         468:    rdata = 32'h00d79463;
         469:    rdata = 32'h0405872a;
         470:    rdata = 32'h46294501;
         471:    rdata = 32'h00044683;
         472:    rdata = 32'h07b3ca81;
         473:    rdata = 32'h851302c5;
         474:    rdata = 32'h0405fd06;
         475:    rdata = 32'hb7fd953e;
         476:    rdata = 32'h0533c319;
         477:    rdata = 32'h40b240a0;
         478:    rdata = 32'h01414422;
         479:    rdata = 32'h07138082;
         480:    rdata = 32'h96630300;
         481:    rdata = 32'h470304e7;
         482:    rdata = 32'h07930014;
         483:    rdata = 32'h10630780;
         484:    rdata = 32'h852204f7;
         485:    rdata = 32'hcd053bd1;
         486:    rdata = 32'h45010409;
         487:    rdata = 32'h06000713;
         488:    rdata = 32'h04000693;
         489:    rdata = 32'h00044783;
         490:    rdata = 32'h7a63d7f9;
         491:    rdata = 32'h879300f7;
         492:    rdata = 32'hf793fa97;
         493:    rdata = 32'h05120ff7;
         494:    rdata = 32'h04058d5d;
         495:    rdata = 32'hf563b7e5;
         496:    rdata = 32'h879300f6;
         497:    rdata = 32'hb7f5fc97;
         498:    rdata = 32'hfd078793;
         499:    rdata = 32'hc537b7dd;
         500:    rdata = 32'h0513dead;
         501:    rdata = 32'hb745eef5;
         502:    rdata = 32'hfdf57793;
         503:    rdata = 32'hfbf78793;
         504:    rdata = 32'h0ff7f793;
         505:    rdata = 32'h77634765;
         506:    rdata = 32'h051300f7;
         507:    rdata = 32'h3513fd05;
         508:    rdata = 32'h808200a5;
         509:    rdata = 32'h80824505;
         510:    rdata = 32'hc150c10c;
         511:    rdata = 32'hf7938082;
         512:    rdata = 32'h410cffc5;
         513:    rdata = 32'h418895be;
         514:    rdata = 32'hf7938082;
         515:    rdata = 32'h410cffc5;
         516:    rdata = 32'hc19095be;
         517:    rdata = 32'h41488082;
         518:    rdata = 32'h25738082;
         519:    rdata = 32'h25f3b000;
         520:    rdata = 32'h8082b800;
         521:    rdata = 32'h00010001;
         522:    rdata = 32'h00010001;
         523:    rdata = 32'h00010001;
         524:    rdata = 32'hf9ed15fd;
         525:    rdata = 32'hc10c8082;
         526:    rdata = 32'h62f38082;
         527:    rdata = 32'h80823004;
         528:    rdata = 32'h300472f3;
         529:    rdata = 32'hc14c8082;
         530:    rdata = 32'ha2f362c1;
         531:    rdata = 32'h80823042;
         532:    rdata = 32'h00052223;
         533:    rdata = 32'hb2f362c1;
         534:    rdata = 32'h80823042;
         535:    rdata = 32'h02b7c50c;
         536:    rdata = 32'ha2f30002;
         537:    rdata = 32'h80823042;
         538:    rdata = 32'h00052423;
         539:    rdata = 32'h000202b7;
         540:    rdata = 32'h3042b2f3;
         541:    rdata = 32'hc54c8082;
         542:    rdata = 32'h000402b7;
         543:    rdata = 32'h3042a2f3;
         544:    rdata = 32'h26238082;
         545:    rdata = 32'h02b70005;
         546:    rdata = 32'hb2f30004;
         547:    rdata = 32'h80823042;
         548:    rdata = 32'h02b7c90c;
         549:    rdata = 32'ha2f30008;
         550:    rdata = 32'h80823042;
         551:    rdata = 32'h00052823;
         552:    rdata = 32'h000802b7;
         553:    rdata = 32'h3042b2f3;
         554:    rdata = 32'h71398082;
         555:    rdata = 32'hde06d036;
         556:    rdata = 32'hda1adc16;
         557:    rdata = 32'hd62ad81e;
         558:    rdata = 32'hd232d42e;
         559:    rdata = 32'hcc3ece3a;
         560:    rdata = 32'hc846ca42;
         561:    rdata = 32'hc476c672;
         562:    rdata = 32'hc07ec27a;
         563:    rdata = 32'h000ff697;
         564:    rdata = 32'h7346a683;
         565:    rdata = 32'h2673ce9d;
         566:    rdata = 32'h42183410;
         567:    rdata = 32'h8b0d4791;
         568:    rdata = 32'h4789e311;
         569:    rdata = 32'h907397b2;
         570:    rdata = 32'h96823417;
         571:    rdata = 32'h52e250f2;
         572:    rdata = 32'h53c25352;
         573:    rdata = 32'h55a25532;
         574:    rdata = 32'h56825612;
         575:    rdata = 32'h47e24772;
         576:    rdata = 32'h48c24852;
         577:    rdata = 32'h4ea24e32;
         578:    rdata = 32'h4f824f12;
         579:    rdata = 32'h00736121;
         580:    rdata = 32'ha0013020;
         581:    rdata = 32'hcc3e7139;
         582:    rdata = 32'hdc16de06;
         583:    rdata = 32'hd81eda1a;
         584:    rdata = 32'hd42ed62a;
         585:    rdata = 32'hd036d232;
         586:    rdata = 32'hca42ce3a;
         587:    rdata = 32'hc672c846;
         588:    rdata = 32'hc27ac476;
         589:    rdata = 32'hf797c07e;
         590:    rdata = 32'ha783000f;
         591:    rdata = 32'h97826ce7;
         592:    rdata = 32'h52e250f2;
         593:    rdata = 32'h53c25352;
         594:    rdata = 32'h55a25532;
         595:    rdata = 32'h56825612;
         596:    rdata = 32'h47e24772;
         597:    rdata = 32'h48c24852;
         598:    rdata = 32'h4ea24e32;
         599:    rdata = 32'h4f824f12;
         600:    rdata = 32'h00736121;
         601:    rdata = 32'h71393020;
         602:    rdata = 32'hde06cc3e;
         603:    rdata = 32'hda1adc16;
         604:    rdata = 32'hd62ad81e;
         605:    rdata = 32'hd232d42e;
         606:    rdata = 32'hce3ad036;
         607:    rdata = 32'hc846ca42;
         608:    rdata = 32'hc476c672;
         609:    rdata = 32'hc07ec27a;
         610:    rdata = 32'h000ff797;
         611:    rdata = 32'h6807a783;
         612:    rdata = 32'h50f29782;
         613:    rdata = 32'h535252e2;
         614:    rdata = 32'h553253c2;
         615:    rdata = 32'h561255a2;
         616:    rdata = 32'h47725682;
         617:    rdata = 32'h485247e2;
         618:    rdata = 32'h4e3248c2;
         619:    rdata = 32'h4f124ea2;
         620:    rdata = 32'h61214f82;
         621:    rdata = 32'h30200073;
         622:    rdata = 32'hcc3e7139;
         623:    rdata = 32'hdc16de06;
         624:    rdata = 32'hd81eda1a;
         625:    rdata = 32'hd42ed62a;
         626:    rdata = 32'hd036d232;
         627:    rdata = 32'hca42ce3a;
         628:    rdata = 32'hc672c846;
         629:    rdata = 32'hc27ac476;
         630:    rdata = 32'hf797c07e;
         631:    rdata = 32'ha783000f;
         632:    rdata = 32'h97826327;
         633:    rdata = 32'h52e250f2;
         634:    rdata = 32'h53c25352;
         635:    rdata = 32'h55a25532;
         636:    rdata = 32'h56825612;
         637:    rdata = 32'h47e24772;
         638:    rdata = 32'h48c24852;
         639:    rdata = 32'h4ea24e32;
         640:    rdata = 32'h4f824f12;
         641:    rdata = 32'h00736121;
         642:    rdata = 32'h71393020;
         643:    rdata = 32'hde06cc3e;
         644:    rdata = 32'hda1adc16;
         645:    rdata = 32'hd62ad81e;
         646:    rdata = 32'hd232d42e;
         647:    rdata = 32'hce3ad036;
         648:    rdata = 32'hc846ca42;
         649:    rdata = 32'hc476c672;
         650:    rdata = 32'hc07ec27a;
         651:    rdata = 32'h000ff797;
         652:    rdata = 32'h5e47a783;
         653:    rdata = 32'h50f29782;
         654:    rdata = 32'h535252e2;
         655:    rdata = 32'h553253c2;
         656:    rdata = 32'h561255a2;
         657:    rdata = 32'h47725682;
         658:    rdata = 32'h485247e2;
         659:    rdata = 32'h4e3248c2;
         660:    rdata = 32'h4f124ea2;
         661:    rdata = 32'h61214f82;
         662:    rdata = 32'h30200073;
         663:    rdata = 32'h8082c10c;
         664:    rdata = 32'h00163613;
         665:    rdata = 32'h000ff517;
         666:    rdata = 32'h5b850513;
         667:    rdata = 32'h1141a8d9;
         668:    rdata = 32'h000ff517;
         669:    rdata = 32'h5ac50513;
         670:    rdata = 32'h20f5c606;
         671:    rdata = 32'h157d40b2;
         672:    rdata = 32'h00a03533;
         673:    rdata = 32'h80820141;
         674:    rdata = 32'h87324108;
         675:    rdata = 32'h862e4685;
         676:    rdata = 32'ha9cd4581;
         677:    rdata = 32'hcc221101;
         678:    rdata = 32'h842ac62e;
         679:    rdata = 32'h3fc1ce06;
         680:    rdata = 32'h463287aa;
         681:    rdata = 32'h46854008;
         682:    rdata = 32'hc3914581;
         683:    rdata = 32'h21d94591;
         684:    rdata = 32'h446240f2;
         685:    rdata = 32'h00a03533;
         686:    rdata = 32'h80826105;
         687:    rdata = 32'h862e4108;
         688:    rdata = 32'h45814685;
         689:    rdata = 32'h4108a9f1;
         690:    rdata = 32'h4705862e;
         691:    rdata = 32'h45a14685;
         692:    rdata = 32'h4108a955;
         693:    rdata = 32'h4701862e;
         694:    rdata = 32'h45a14685;
         695:    rdata = 32'h4108a165;
         696:    rdata = 32'h862e1141;
         697:    rdata = 32'h45b14685;
         698:    rdata = 32'h2169c606;
         699:    rdata = 32'h353340b2;
         700:    rdata = 32'h014100a0;
         701:    rdata = 32'h41088082;
         702:    rdata = 32'h4701862e;
         703:    rdata = 32'h45b14685;
         704:    rdata = 32'h4108a151;
         705:    rdata = 32'h4705862e;
         706:    rdata = 32'h45c14685;
         707:    rdata = 32'h4108a9a5;
         708:    rdata = 32'h4701862e;
         709:    rdata = 32'h45c14685;
         710:    rdata = 32'h4108a1b5;
         711:    rdata = 32'h862e1141;
         712:    rdata = 32'h45d14685;
         713:    rdata = 32'h21b9c606;
         714:    rdata = 32'h353340b2;
         715:    rdata = 32'h014100a0;
         716:    rdata = 32'h41088082;
         717:    rdata = 32'h4701862e;
         718:    rdata = 32'h45d14685;
         719:    rdata = 32'hc10ca1a1;
         720:    rdata = 32'h47bd8082;
         721:    rdata = 32'h87324108;
         722:    rdata = 32'h00b7e863;
         723:    rdata = 32'hf6130586;
         724:    rdata = 32'h468d0fe5;
         725:    rdata = 32'ha13d4581;
         726:    rdata = 32'h058615c1;
         727:    rdata = 32'h0fe5f613;
         728:    rdata = 32'h4591468d;
         729:    rdata = 32'h1141bfcd;
         730:    rdata = 32'h47bdc606;
         731:    rdata = 32'he6634108;
         732:    rdata = 32'h961302b7;
         733:    rdata = 32'h468d0015;
         734:    rdata = 32'h0fe67613;
         735:    rdata = 32'h2edd4581;
         736:    rdata = 32'h470587aa;
         737:    rdata = 32'h87634505;
         738:    rdata = 32'h470900e7;
         739:    rdata = 32'h93634501;
         740:    rdata = 32'h450900e7;
         741:    rdata = 32'h014140b2;
         742:    rdata = 32'h86138082;
         743:    rdata = 32'h0606ff05;
         744:    rdata = 32'h7613468d;
         745:    rdata = 32'h45910fe6;
         746:    rdata = 32'hc10cbfd9;
         747:    rdata = 32'h11418082;
         748:    rdata = 32'h45e54609;
         749:    rdata = 32'h000ff517;
         750:    rdata = 32'h46850513;
         751:    rdata = 32'h3751c606;
         752:    rdata = 32'h45ed4609;
         753:    rdata = 32'h000ff517;
         754:    rdata = 32'h45850513;
         755:    rdata = 32'h46093f9d;
         756:    rdata = 32'hf51745f1;
         757:    rdata = 32'h0513000f;
         758:    rdata = 32'h37a544a5;
         759:    rdata = 32'h460940b2;
         760:    rdata = 32'hf51745f5;
         761:    rdata = 32'h0513000f;
         762:    rdata = 32'h014143a5;
         763:    rdata = 32'h4108bf99;
         764:    rdata = 32'h4685872e;
         765:    rdata = 32'h45814601;
         766:    rdata = 32'h4108a671;
         767:    rdata = 32'h4685872e;
         768:    rdata = 32'h45814605;
         769:    rdata = 32'h4108a641;
         770:    rdata = 32'h4685872e;
         771:    rdata = 32'h45814609;
         772:    rdata = 32'h4108ae95;
         773:    rdata = 32'h0693872e;
         774:    rdata = 32'h46010ff0;
         775:    rdata = 32'ha69d45c1;
         776:    rdata = 32'h47014108;
         777:    rdata = 32'h46014685;
         778:    rdata = 32'haea945d1;
         779:    rdata = 32'h11414108;
         780:    rdata = 32'h46014685;
         781:    rdata = 32'hc60645e1;
         782:    rdata = 32'h40b22e35;
         783:    rdata = 32'h00a03533;
         784:    rdata = 32'h80820141;
         785:    rdata = 32'h47014108;
         786:    rdata = 32'h46014685;
         787:    rdata = 32'hae1d45e1;
         788:    rdata = 32'hc4221141;
         789:    rdata = 32'h842ac606;
         790:    rdata = 32'h400837f5;
         791:    rdata = 32'h40b24422;
         792:    rdata = 32'h46854705;
         793:    rdata = 32'h45d14601;
         794:    rdata = 32'hae290141;
         795:    rdata = 32'h872e4108;
         796:    rdata = 32'h0ff00693;
         797:    rdata = 32'h45a14601;
         798:    rdata = 32'h4108a631;
         799:    rdata = 32'h06931141;
         800:    rdata = 32'h46010ff0;
         801:    rdata = 32'hc60645b1;
         802:    rdata = 32'h40b224f5;
         803:    rdata = 32'h0ff57513;
         804:    rdata = 32'h80820141;
         805:    rdata = 32'h11414108;
         806:    rdata = 32'h46054685;
         807:    rdata = 32'hc6064591;
         808:    rdata = 32'h40b22cd1;
         809:    rdata = 32'h00a03533;
         810:    rdata = 32'h80820141;
         811:    rdata = 32'h45811141;
         812:    rdata = 32'hc606c422;
         813:    rdata = 32'h3f5d842a;
         814:    rdata = 32'h3fe98522;
         815:    rdata = 32'h8522fd75;
         816:    rdata = 32'h40b24422;
         817:    rdata = 32'hbf550141;
         818:    rdata = 32'h11414108;
         819:    rdata = 32'h46094685;
         820:    rdata = 32'hc6064591;
         821:    rdata = 32'h40b22445;
         822:    rdata = 32'h00a03533;
         823:    rdata = 32'h80820141;
         824:    rdata = 32'hc4221141;
         825:    rdata = 32'h842ac606;
         826:    rdata = 32'h85223751;
         827:    rdata = 32'hfd753ff1;
         828:    rdata = 32'h44228522;
         829:    rdata = 32'h014140b2;
         830:    rdata = 32'h1101b749;
         831:    rdata = 32'hca26cc22;
         832:    rdata = 32'hc64ec84a;
         833:    rdata = 32'h84aace06;
         834:    rdata = 32'h89b2892e;
         835:    rdata = 32'h5d634401;
         836:    rdata = 32'h85260134;
         837:    rdata = 32'hfd753f55;
         838:    rdata = 32'h008907b3;
         839:    rdata = 32'h0007c583;
         840:    rdata = 32'h04058526;
         841:    rdata = 32'hb7e537a1;
         842:    rdata = 32'h446240f2;
         843:    rdata = 32'h494244d2;
         844:    rdata = 32'h610549b2;
         845:    rdata = 32'h41088082;
         846:    rdata = 32'h46851141;
         847:    rdata = 32'h4591460d;
         848:    rdata = 32'h2c0dc606;
         849:    rdata = 32'h353340b2;
         850:    rdata = 32'h014100a0;
         851:    rdata = 32'h11418082;
         852:    rdata = 32'hc606c422;
         853:    rdata = 32'h8522842a;
         854:    rdata = 32'hdd753ff9;
         855:    rdata = 32'h3f1d8522;
         856:    rdata = 32'h8522e501;
         857:    rdata = 32'hbfdd3f19;
         858:    rdata = 32'h442240b2;
         859:    rdata = 32'h80820141;
         860:    rdata = 32'hc4221141;
         861:    rdata = 32'h842ac606;
         862:    rdata = 32'h85223749;
         863:    rdata = 32'h40b24422;
         864:    rdata = 32'hb7f10141;
         865:    rdata = 32'h8082c10c;
         866:    rdata = 32'hc4221141;
         867:    rdata = 32'h4108842a;
         868:    rdata = 32'h06934731;
         869:    rdata = 32'h46010ff0;
         870:    rdata = 32'hc60645c1;
         871:    rdata = 32'h460922e5;
         872:    rdata = 32'hf51745fd;
         873:    rdata = 32'h0513000f;
         874:    rdata = 32'h3b6127a5;
         875:    rdata = 32'h45f94609;
         876:    rdata = 32'h000ff517;
         877:    rdata = 32'h26c50513;
         878:    rdata = 32'h40083369;
         879:    rdata = 32'h40b24422;
         880:    rdata = 32'h46854705;
         881:    rdata = 32'h45814601;
         882:    rdata = 32'haa6d0141;
         883:    rdata = 32'h11414108;
         884:    rdata = 32'h46014685;
         885:    rdata = 32'hc6064591;
         886:    rdata = 32'h40b22a71;
         887:    rdata = 32'h00a03533;
         888:    rdata = 32'h80820141;
         889:    rdata = 32'h11414108;
         890:    rdata = 32'h0ff00693;
         891:    rdata = 32'h45b14601;
         892:    rdata = 32'h2249c606;
         893:    rdata = 32'h751340b2;
         894:    rdata = 32'h01410ff5;
         895:    rdata = 32'h11418082;
         896:    rdata = 32'hc606c422;
         897:    rdata = 32'h8522842a;
         898:    rdata = 32'hdd7537d1;
         899:    rdata = 32'h44228522;
         900:    rdata = 32'h014140b2;
         901:    rdata = 32'h1101bfc1;
         902:    rdata = 32'hca26cc22;
         903:    rdata = 32'hc64ec84a;
         904:    rdata = 32'hc05ac256;
         905:    rdata = 32'hc452ce06;
         906:    rdata = 32'h892e84aa;
         907:    rdata = 32'h440189b2;
         908:    rdata = 32'h4b214aa9;
         909:    rdata = 32'h03345f63;
         910:    rdata = 32'h0a338526;
         911:    rdata = 32'h37c10089;
         912:    rdata = 32'h00aa0023;
         913:    rdata = 32'h01551f63;
         914:    rdata = 32'h000a0023;
         915:    rdata = 32'h40f24501;
         916:    rdata = 32'h44d24462;
         917:    rdata = 32'h49b24942;
         918:    rdata = 32'h4a924a22;
         919:    rdata = 32'h61054b02;
         920:    rdata = 32'h14638082;
         921:    rdata = 32'hc4010165;
         922:    rdata = 32'h04051479;
         923:    rdata = 32'h547db7e1;
         924:    rdata = 32'h4505bfed;
         925:    rdata = 32'h4108bfe9;
         926:    rdata = 32'h46851141;
         927:    rdata = 32'h45914605;
         928:    rdata = 32'h28cdc606;
         929:    rdata = 32'h353340b2;
         930:    rdata = 32'h014100a0;
         931:    rdata = 32'h41088082;
         932:    rdata = 32'h0693872e;
         933:    rdata = 32'h46010ff0;
         934:    rdata = 32'ha0ed45a1;
         935:    rdata = 32'hcc221101;
         936:    rdata = 32'h842ace06;
         937:    rdata = 32'hc62e8522;
         938:    rdata = 32'h45b237f9;
         939:    rdata = 32'h8522fd65;
         940:    rdata = 32'h40f24462;
         941:    rdata = 32'hbfe16105;
         942:    rdata = 32'hc4221141;
         943:    rdata = 32'hc606c226;
         944:    rdata = 32'h842e84aa;
         945:    rdata = 32'h00044583;
         946:    rdata = 32'h8526c589;
         947:    rdata = 32'h37f90405;
         948:    rdata = 32'h40b2bfd5;
         949:    rdata = 32'h44924422;
         950:    rdata = 32'h80820141;
         951:    rdata = 32'h47014108;
         952:    rdata = 32'h46014685;
         953:    rdata = 32'ha87945d1;
         954:    rdata = 32'h11414108;
         955:    rdata = 32'h46014685;
         956:    rdata = 32'hc60645e1;
         957:    rdata = 32'h40b22041;
         958:    rdata = 32'h00a03533;
         959:    rdata = 32'h80820141;
         960:    rdata = 32'h47014108;
         961:    rdata = 32'h46014685;
         962:    rdata = 32'ha8ad45e1;
         963:    rdata = 32'hc4221141;
         964:    rdata = 32'h842ac606;
         965:    rdata = 32'h400837f5;
         966:    rdata = 32'h40b24422;
         967:    rdata = 32'h46854705;
         968:    rdata = 32'h45d14601;
         969:    rdata = 32'ha8b90141;
         970:    rdata = 32'h47014108;
         971:    rdata = 32'h46054685;
         972:    rdata = 32'ha88945d1;
         973:    rdata = 32'h11414108;
         974:    rdata = 32'h46054685;
         975:    rdata = 32'hc60645e1;
         976:    rdata = 32'h40b22815;
         977:    rdata = 32'h00a03533;
         978:    rdata = 32'h80820141;
         979:    rdata = 32'h47014108;
         980:    rdata = 32'h46054685;
         981:    rdata = 32'ha03d45e1;
         982:    rdata = 32'hc4221141;
         983:    rdata = 32'h842ac606;
         984:    rdata = 32'h400837f5;
         985:    rdata = 32'h40b24422;
         986:    rdata = 32'h46854705;
         987:    rdata = 32'h45d14605;
         988:    rdata = 32'ha8090141;
         989:    rdata = 32'h952e99f1;
         990:    rdata = 32'hd7b3411c;
         991:    rdata = 32'hf53300c7;
         992:    rdata = 32'h808200d7;
         993:    rdata = 32'h952e99f1;
         994:    rdata = 32'h97b3410c;
         995:    rdata = 32'hc79300c6;
         996:    rdata = 32'h8ef9fff7;
         997:    rdata = 32'h96b38fed;
         998:    rdata = 32'h8edd00c6;
         999:    rdata = 32'h8082c114;
        1000:    rdata = 32'h952e99f1;
        1001:    rdata = 32'h96b3411c;
        1002:    rdata = 32'h8ebd00c6;
        1003:    rdata = 32'h8082c114;
        1004:    rdata = 32'hf5171101;
        1005:    rdata = 32'h0513000f;
        1006:    rdata = 32'hce0606e5;
        1007:    rdata = 32'hf5173ecd;
        1008:    rdata = 32'h0513000f;
        1009:    rdata = 32'h33c90665;
        1010:    rdata = 32'h00000597;
        1011:    rdata = 32'h17058593;
        1012:    rdata = 32'h000ff517;
        1013:    rdata = 32'h04450513;
        1014:    rdata = 32'hc84ff0ef;
        1015:    rdata = 32'h850a45e9;
        1016:    rdata = 32'haeaff0ef;
        1017:    rdata = 32'hf0ef850a;
        1018:    rdata = 32'h45ddaf6f;
        1019:    rdata = 32'h000ff517;
        1020:    rdata = 32'h02c50513;
        1021:    rdata = 32'haa1ff0ef;
        1022:    rdata = 32'h0597c539;
        1023:    rdata = 32'h85930000;
        1024:    rdata = 32'hf51715a5;
        1025:    rdata = 32'h0513000f;
        1026:    rdata = 32'hf0ef0125;
        1027:    rdata = 32'h62c1c52f;
        1028:    rdata = 32'h305292f3;
        1029:    rdata = 32'h00000597;
        1030:    rdata = 32'h1e458593;
        1031:    rdata = 32'h000ff517;
        1032:    rdata = 32'hff850513;
        1033:    rdata = 32'hc38ff0ef;
        1034:    rdata = 32'h000ff517;
        1035:    rdata = 32'hfec50513;
        1036:    rdata = 32'hc70ff0ef;
        1037:    rdata = 32'hf0ef850a;
        1038:    rdata = 32'hf06fb9ef;
        1039:    rdata = 32'h40f20460;
        1040:    rdata = 32'h61054501;
        1041:    rdata = 32'h00288082;
        1042:    rdata = 32'h94cff0ef;
        1043:    rdata = 32'hf51745e1;
        1044:    rdata = 32'h0513000f;
        1045:    rdata = 32'hf0effca5;
        1046:    rdata = 32'hc525a3ff;
        1047:    rdata = 32'h00000597;
        1048:    rdata = 32'h11058593;
        1049:    rdata = 32'h000ff517;
        1050:    rdata = 32'hfb050513;
        1051:    rdata = 32'hbf0ff0ef;
        1052:    rdata = 32'hf0ef0028;
        1053:    rdata = 32'hc22a9a8f;
        1054:    rdata = 32'h0597c51d;
        1055:    rdata = 32'h85930000;
        1056:    rdata = 32'hf5171125;
        1057:    rdata = 32'h0513000f;
        1058:    rdata = 32'hf0eff925;
        1059:    rdata = 32'h004cbd2f;
        1060:    rdata = 32'hbeaff0ef;
        1061:    rdata = 32'h00000597;
        1062:    rdata = 32'h0bc58593;
        1063:    rdata = 32'hbc0ff0ef;
        1064:    rdata = 32'hf0ef850a;
        1065:    rdata = 32'h0597af8f;
        1066:    rdata = 32'h85930000;
        1067:    rdata = 32'hf5171365;
        1068:    rdata = 32'h0513000f;
        1069:    rdata = 32'hf0eff665;
        1070:    rdata = 32'h850aba6f;
        1071:    rdata = 32'ha64ff0ef;
        1072:    rdata = 32'h0597b7b9;
        1073:    rdata = 32'h85930000;
        1074:    rdata = 32'hf5170fe5;
        1075:    rdata = 32'h0513000f;
        1076:    rdata = 32'hf0eff4a5;
        1077:    rdata = 32'h0028b8af;
        1078:    rdata = 32'h8c2ff0ef;
        1079:    rdata = 32'h17b7b7e9;
        1080:    rdata = 32'hf7170100;
        1081:    rdata = 32'h2b23000f;
        1082:    rdata = 32'h8082f2f7;
        1083:    rdata = 32'h010007b7;
        1084:    rdata = 32'h000ff717;
        1085:    rdata = 32'hf2f72623;
        1086:    rdata = 32'h37b78082;
        1087:    rdata = 32'hf7170100;
        1088:    rdata = 32'h2123000f;
        1089:    rdata = 32'h8082f2f7;
        1090:    rdata = 32'h010027b7;
        1091:    rdata = 32'h000ff717;
        1092:    rdata = 32'hf0f72c23;
        1093:    rdata = 32'h00008082;
        1094:    rdata = 32'h00000000;
        1095:    rdata = 32'h00000000;
        1096:    rdata = 32'h00000000;
        1097:    rdata = 32'h00000000;
        1098:    rdata = 32'h000010de;
        1099:    rdata = 32'h000010ec;
        1100:    rdata = 32'h000010fa;
        1101:    rdata = 32'h00001108;
        1102:    rdata = 32'h4f464e49;
        1103:    rdata = 32'h6f62203a;
        1104:    rdata = 32'h6f6c746f;
        1105:    rdata = 32'h72656461;
        1106:    rdata = 32'h61747320;
        1107:    rdata = 32'h64657472;
        1108:    rdata = 32'h0000000a;
        1109:    rdata = 32'h4f464e49;
        1110:    rdata = 32'h6f63203a;
        1111:    rdata = 32'h6f6c6564;
        1112:    rdata = 32'h73206461;
        1113:    rdata = 32'h7070696b;
        1114:    rdata = 32'h000a6465;
        1115:    rdata = 32'h4f464e49;
        1116:    rdata = 32'h6f63203a;
        1117:    rdata = 32'h6f6c6564;
        1118:    rdata = 32'h73206461;
        1119:    rdata = 32'h6372756f;
        1120:    rdata = 32'h75203a65;
        1121:    rdata = 32'h0a747261;
        1122:    rdata = 32'h00000000;
        1123:    rdata = 32'h4f525245;
        1124:    rdata = 32'h63203a52;
        1125:    rdata = 32'h6c65646f;
        1126:    rdata = 32'h2064616f;
        1127:    rdata = 32'h656d6974;
        1128:    rdata = 32'h2074756f;
        1129:    rdata = 32'h7563636f;
        1130:    rdata = 32'h64657272;
        1131:    rdata = 32'h6572202e;
        1132:    rdata = 32'h76696563;
        1133:    rdata = 32'h62206465;
        1134:    rdata = 32'h73657479;
        1135:    rdata = 32'h0000203a;
        1136:    rdata = 32'h4f464e49;
        1137:    rdata = 32'h6f63203a;
        1138:    rdata = 32'h6f6c6564;
        1139:    rdata = 32'h73206461;
        1140:    rdata = 32'h6372756f;
        1141:    rdata = 32'h73203a65;
        1142:    rdata = 32'h000a6970;
        1143:    rdata = 32'h4f464e49;
        1144:    rdata = 32'h6f63203a;
        1145:    rdata = 32'h6f6c6564;
        1146:    rdata = 32'h66206461;
        1147:    rdata = 32'h73696e69;
        1148:    rdata = 32'h0a646568;
        1149:    rdata = 32'h00000000;
        1150:    rdata = 32'h4f464e49;
        1151:    rdata = 32'h6f62203a;
        1152:    rdata = 32'h6f6c746f;
        1153:    rdata = 32'h72656461;
        1154:    rdata = 32'h6e696620;
        1155:    rdata = 32'h65687369;
        1156:    rdata = 32'h00000a64;
        1157:    rdata = 32'h6f636e69;
        1158:    rdata = 32'h63657272;
        1159:    rdata = 32'h61762074;
        1160:    rdata = 32'h2e65756c;
        1161:    rdata = 32'h79727420;
        1162:    rdata = 32'h61676120;
        1163:    rdata = 32'h000a6e69;
        default: rdata = 32'h00000000;
    endcase
end
endmodule
