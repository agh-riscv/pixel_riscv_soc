/**
 * Copyright (C) 2020  AGH University of Science and Technology
 *
 * This program is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with this program.  If not, see <https://www.gnu.org/licenses/>.
 */

module boot_mem (
    output logic [31:0] rdata,
    input logic [31:0] addr
);

/**
 * Module internal logic
 */

always_comb begin
    case (addr[13:2])
           0:    rdata = 32'h08c0006f;
           1:    rdata = 32'h0880006f;
           2:    rdata = 32'h0840006f;
           3:    rdata = 32'h0800006f;
           4:    rdata = 32'h07c0006f;
           5:    rdata = 32'h0780006f;
           6:    rdata = 32'h0740006f;
           7:    rdata = 32'h0700006f;
           8:    rdata = 32'h06c0006f;
           9:    rdata = 32'h0680006f;
          10:    rdata = 32'h0640006f;
          11:    rdata = 32'h0600006f;
          12:    rdata = 32'h05c0006f;
          13:    rdata = 32'h0580006f;
          14:    rdata = 32'h0540006f;
          15:    rdata = 32'h0500006f;
          16:    rdata = 32'h04c0006f;
          17:    rdata = 32'h0480006f;
          18:    rdata = 32'h0440006f;
          19:    rdata = 32'h0400006f;
          20:    rdata = 32'h03c0006f;
          21:    rdata = 32'h0380006f;
          22:    rdata = 32'h0340006f;
          23:    rdata = 32'h0300006f;
          24:    rdata = 32'h02c0006f;
          25:    rdata = 32'h0280006f;
          26:    rdata = 32'h0240006f;
          27:    rdata = 32'h0200006f;
          28:    rdata = 32'h01c0006f;
          29:    rdata = 32'h0180006f;
          30:    rdata = 32'h0140006f;
          31:    rdata = 32'h0100006f;
          32:    rdata = 32'h0100006f;
          33:    rdata = 32'h0080006f;
          34:    rdata = 32'h0040006f;
          35:    rdata = 32'h0000006f;
          36:    rdata = 32'h00000093;
          37:    rdata = 32'h00000113;
          38:    rdata = 32'h00000193;
          39:    rdata = 32'h00000213;
          40:    rdata = 32'h00000293;
          41:    rdata = 32'h00000313;
          42:    rdata = 32'h00000393;
          43:    rdata = 32'h00000413;
          44:    rdata = 32'h00000493;
          45:    rdata = 32'h00000513;
          46:    rdata = 32'h00000593;
          47:    rdata = 32'h00000613;
          48:    rdata = 32'h00000693;
          49:    rdata = 32'h00000713;
          50:    rdata = 32'h00000793;
          51:    rdata = 32'h00000813;
          52:    rdata = 32'h00000893;
          53:    rdata = 32'h00000913;
          54:    rdata = 32'h00000993;
          55:    rdata = 32'h00000a13;
          56:    rdata = 32'h00000a93;
          57:    rdata = 32'h00000b13;
          58:    rdata = 32'h00000b93;
          59:    rdata = 32'h00000c13;
          60:    rdata = 32'h00000c93;
          61:    rdata = 32'h00000d13;
          62:    rdata = 32'h00000d93;
          63:    rdata = 32'h00000e13;
          64:    rdata = 32'h00000e93;
          65:    rdata = 32'h00000f13;
          66:    rdata = 32'h00000f93;
          67:    rdata = 32'h00104117;
          68:    rdata = 32'hef410113;
          69:    rdata = 32'h00100297;
          70:    rdata = 32'heec28293;
          71:    rdata = 32'h00100317;
          72:    rdata = 32'hf4830313;
          73:    rdata = 32'h0062d863;
          74:    rdata = 32'h0002a023;
          75:    rdata = 32'h00428293;
          76:    rdata = 32'hfe535ce3;
          77:    rdata = 32'h00001297;
          78:    rdata = 32'hc3028293;
          79:    rdata = 32'h00100317;
          80:    rdata = 32'hec430313;
          81:    rdata = 32'h00100397;
          82:    rdata = 32'hebc38393;
          83:    rdata = 32'h00735c63;
          84:    rdata = 32'h0002ae03;
          85:    rdata = 32'h01c32023;
          86:    rdata = 32'h00428293;
          87:    rdata = 32'h00430313;
          88:    rdata = 32'hfe7348e3;
          89:    rdata = 32'h00001297;
          90:    rdata = 32'hb0428293;
          91:    rdata = 32'h00001317;
          92:    rdata = 32'hb0c30313;
          93:    rdata = 32'h0062da63;
          94:    rdata = 32'h0002a783;
          95:    rdata = 32'h000780e7;
          96:    rdata = 32'h00428293;
          97:    rdata = 32'hfe62cae3;
          98:    rdata = 32'h00000513;
          99:    rdata = 32'h00000593;
         100:    rdata = 32'h19b000ef;
         101:    rdata = 32'h45857179;
         102:    rdata = 32'h00100517;
         103:    rdata = 32'he9850513;
         104:    rdata = 32'hd422d606;
         105:    rdata = 32'hce4ed04a;
         106:    rdata = 32'hd226cc52;
         107:    rdata = 32'h029000ef;
         108:    rdata = 32'h0517458d;
         109:    rdata = 32'h05130010;
         110:    rdata = 32'h00efe7e5;
         111:    rdata = 32'h440103d0;
         112:    rdata = 32'h00100917;
         113:    rdata = 32'he9c90913;
         114:    rdata = 32'h00100997;
         115:    rdata = 32'he6898993;
         116:    rdata = 32'h854a4a11;
         117:    rdata = 32'h74632365;
         118:    rdata = 32'h448102a4;
         119:    rdata = 32'h00ef854e;
         120:    rdata = 32'h007c0210;
         121:    rdata = 32'h802397a6;
         122:    rdata = 32'h048500a7;
         123:    rdata = 32'hff4498e3;
         124:    rdata = 32'h85a244b2;
         125:    rdata = 32'h2bbd854a;
         126:    rdata = 32'h0411c104;
         127:    rdata = 32'h50b2bfd9;
         128:    rdata = 32'h54925422;
         129:    rdata = 32'h49f25902;
         130:    rdata = 32'h61454a62;
         131:    rdata = 32'h71398082;
         132:    rdata = 32'h0517da26;
         133:    rdata = 32'h05130010;
         134:    rdata = 32'hd4b7dee5;
         135:    rdata = 32'hdc223b9a;
         136:    rdata = 32'hd452d84a;
         137:    rdata = 32'hd05ad256;
         138:    rdata = 32'hde06ce5e;
         139:    rdata = 32'h8493d64e;
         140:    rdata = 32'h23b9a004;
         141:    rdata = 32'hb53394aa;
         142:    rdata = 32'h043300a4;
         143:    rdata = 32'h490100b5;
         144:    rdata = 32'h00100a97;
         145:    rdata = 32'he1ca8a93;
         146:    rdata = 32'h00100a17;
         147:    rdata = 32'hdfca0a13;
         148:    rdata = 32'h00100b17;
         149:    rdata = 32'hdb0b0b13;
         150:    rdata = 32'h85564b91;
         151:    rdata = 32'h71632305;
         152:    rdata = 32'h498106a9;
         153:    rdata = 32'h00ef8552;
         154:    rdata = 32'he9090b10;
         155:    rdata = 32'h2b09855a;
         156:    rdata = 32'hfe85eae3;
         157:    rdata = 32'h00b41463;
         158:    rdata = 32'hfe9566e3;
         159:    rdata = 32'h00ef8552;
         160:    rdata = 32'hc11d0990;
         161:    rdata = 32'h00ef8552;
         162:    rdata = 32'h007c0990;
         163:    rdata = 32'h802397ce;
         164:    rdata = 32'h098500a7;
         165:    rdata = 32'hfd7998e3;
         166:    rdata = 32'h85ca49b2;
         167:    rdata = 32'h29d98556;
         168:    rdata = 32'h01352023;
         169:    rdata = 32'hbf550911;
         170:    rdata = 32'h50f2557d;
         171:    rdata = 32'h54d25462;
         172:    rdata = 32'h59b25942;
         173:    rdata = 32'h5a925a22;
         174:    rdata = 32'h4bf25b02;
         175:    rdata = 32'h80826121;
         176:    rdata = 32'hb7e54501;
         177:    rdata = 32'h05131141;
         178:    rdata = 32'hc6060fa0;
         179:    rdata = 32'h458520f9;
         180:    rdata = 32'h00100517;
         181:    rdata = 32'hd3c50513;
         182:    rdata = 32'h051325c1;
         183:    rdata = 32'h28750fa0;
         184:    rdata = 32'h00100517;
         185:    rdata = 32'hd2c50513;
         186:    rdata = 32'h257d4581;
         187:    rdata = 32'h051340b2;
         188:    rdata = 32'h01410fa0;
         189:    rdata = 32'h1141a05d;
         190:    rdata = 32'h0fa00513;
         191:    rdata = 32'h2871c606;
         192:    rdata = 32'h05174585;
         193:    rdata = 32'h05130010;
         194:    rdata = 32'h2579d0a5;
         195:    rdata = 32'h0fa00513;
         196:    rdata = 32'h45812069;
         197:    rdata = 32'h00100517;
         198:    rdata = 32'hcf850513;
         199:    rdata = 32'h05132db5;
         200:    rdata = 32'h28a50fa0;
         201:    rdata = 32'h05174585;
         202:    rdata = 32'h05130010;
         203:    rdata = 32'h25adce65;
         204:    rdata = 32'h0fa00513;
         205:    rdata = 32'h4581209d;
         206:    rdata = 32'h00100517;
         207:    rdata = 32'hcd450513;
         208:    rdata = 32'h05132da1;
         209:    rdata = 32'h28910fa0;
         210:    rdata = 32'h051340b2;
         211:    rdata = 32'h01410fa0;
         212:    rdata = 32'h1141a0a9;
         213:    rdata = 32'h0fa00513;
         214:    rdata = 32'hc606c422;
         215:    rdata = 32'h00100417;
         216:    rdata = 32'hcb040413;
         217:    rdata = 32'h4585281d;
         218:    rdata = 32'h253d8522;
         219:    rdata = 32'h0fa00513;
         220:    rdata = 32'h8522202d;
         221:    rdata = 32'h250d4581;
         222:    rdata = 32'h0fa00513;
         223:    rdata = 32'hb7e52839;
         224:    rdata = 32'h05131141;
         225:    rdata = 32'hc6060fa0;
         226:    rdata = 32'h40b22809;
         227:    rdata = 32'h05174585;
         228:    rdata = 32'h05130010;
         229:    rdata = 32'h0141c7e5;
         230:    rdata = 32'h6785a501;
         231:    rdata = 32'h38878793;
         232:    rdata = 32'h02f505b3;
         233:    rdata = 32'h00100517;
         234:    rdata = 32'hc5c50513;
         235:    rdata = 32'h4595aef9;
         236:    rdata = 32'h02b505b3;
         237:    rdata = 32'h00100517;
         238:    rdata = 32'hc4c50513;
         239:    rdata = 32'h1141a6f9;
         240:    rdata = 32'h0613c422;
         241:    rdata = 32'h842a0640;
         242:    rdata = 32'h00100517;
         243:    rdata = 32'hc7c50513;
         244:    rdata = 32'h257dc606;
         245:    rdata = 32'h852240b2;
         246:    rdata = 32'h01414422;
         247:    rdata = 32'h11418082;
         248:    rdata = 32'h842ac422;
         249:    rdata = 32'h00100517;
         250:    rdata = 32'hc6050513;
         251:    rdata = 32'h2711c606;
         252:    rdata = 32'h852240b2;
         253:    rdata = 32'h01414422;
         254:    rdata = 32'h11418082;
         255:    rdata = 32'h842ac422;
         256:    rdata = 32'h00100517;
         257:    rdata = 32'hc4450513;
         258:    rdata = 32'h25e5c606;
         259:    rdata = 32'h852240b2;
         260:    rdata = 32'h01414422;
         261:    rdata = 32'h418c8082;
         262:    rdata = 32'hcc221101;
         263:    rdata = 32'h0048842a;
         264:    rdata = 32'h2c19ce06;
         265:    rdata = 32'h0517004c;
         266:    rdata = 32'h05130010;
         267:    rdata = 32'h25d1c1e5;
         268:    rdata = 32'h852240f2;
         269:    rdata = 32'h61054462;
         270:    rdata = 32'h71758082;
         271:    rdata = 32'hc326c522;
         272:    rdata = 32'hdecec14a;
         273:    rdata = 32'hc706dcd2;
         274:    rdata = 32'h892e84aa;
         275:    rdata = 32'h00100417;
         276:    rdata = 32'hbf840413;
         277:    rdata = 32'h00001a17;
         278:    rdata = 32'h8f0a0a13;
         279:    rdata = 32'h00001997;
         280:    rdata = 32'h8ec98993;
         281:    rdata = 32'h852285ca;
         282:    rdata = 32'h85d22569;
         283:    rdata = 32'h25518522;
         284:    rdata = 32'h8526006c;
         285:    rdata = 32'h006837a9;
         286:    rdata = 32'he5092409;
         287:    rdata = 32'h852285ce;
         288:    rdata = 32'hb7cd2d8d;
         289:    rdata = 32'h242d0068;
         290:    rdata = 32'h442a40ba;
         291:    rdata = 32'h490a449a;
         292:    rdata = 32'h5a6659f6;
         293:    rdata = 32'h80826149;
         294:    rdata = 32'h03000713;
         295:    rdata = 32'h00054783;
         296:    rdata = 32'h00e79463;
         297:    rdata = 32'hbfdd0505;
         298:    rdata = 32'h157de391;
         299:    rdata = 32'h47038082;
         300:    rdata = 32'h07930005;
         301:    rdata = 32'h136302d0;
         302:    rdata = 32'h050500f7;
         303:    rdata = 32'h47834725;
         304:    rdata = 32'h87930005;
         305:    rdata = 32'hf793fd07;
         306:    rdata = 32'h68630ff7;
         307:    rdata = 32'h478300f7;
         308:    rdata = 32'h05050015;
         309:    rdata = 32'h4505f7ed;
         310:    rdata = 32'h45018082;
         311:    rdata = 32'h05098082;
         312:    rdata = 32'h461546a5;
         313:    rdata = 32'h00054783;
         314:    rdata = 32'hfd078713;
         315:    rdata = 32'h0ff77713;
         316:    rdata = 32'h00e6fa63;
         317:    rdata = 32'hfdf7f793;
         318:    rdata = 32'hfbf78793;
         319:    rdata = 32'h0ff7f793;
         320:    rdata = 32'h00f66863;
         321:    rdata = 32'h00154783;
         322:    rdata = 32'hffe90505;
         323:    rdata = 32'h80824505;
         324:    rdata = 32'h80824501;
         325:    rdata = 32'hc70387aa;
         326:    rdata = 32'h05850005;
         327:    rdata = 32'h8fa30785;
         328:    rdata = 32'hfb75fee7;
         329:    rdata = 32'h87aa8082;
         330:    rdata = 32'h0007c683;
         331:    rdata = 32'h0785873e;
         332:    rdata = 32'hc783fee5;
         333:    rdata = 32'h05850005;
         334:    rdata = 32'h0fa30705;
         335:    rdata = 32'hfbf5fef7;
         336:    rdata = 32'h47838082;
         337:    rdata = 32'hc7030005;
         338:    rdata = 32'h87630005;
         339:    rdata = 32'h557d00e7;
         340:    rdata = 32'h00e7e963;
         341:    rdata = 32'h80824505;
         342:    rdata = 32'h0505c781;
         343:    rdata = 32'hb7d50585;
         344:    rdata = 32'h80824501;
         345:    rdata = 32'h450187aa;
         346:    rdata = 32'h00a78733;
         347:    rdata = 32'h00074703;
         348:    rdata = 32'h0505c319;
         349:    rdata = 32'h8082bfd5;
         350:    rdata = 32'h0c634789;
         351:    rdata = 32'h479102f6;
         352:    rdata = 32'h02f60d63;
         353:    rdata = 32'h47814705;
         354:    rdata = 32'h00e61463;
         355:    rdata = 32'h06400793;
         356:    rdata = 32'hcb8d4629;
         357:    rdata = 32'h02f5d733;
         358:    rdata = 32'h76930505;
         359:    rdata = 32'h86b30ff7;
         360:    rdata = 32'h071302f6;
         361:    rdata = 32'h0fa30307;
         362:    rdata = 32'hd7b3fee5;
         363:    rdata = 32'h8d9502c7;
         364:    rdata = 32'h6789b7cd;
         365:    rdata = 32'h71078793;
         366:    rdata = 32'hd7b7bfe1;
         367:    rdata = 32'h87933b9a;
         368:    rdata = 32'hb7f9a007;
         369:    rdata = 32'h00050023;
         370:    rdata = 32'h46058082;
         371:    rdata = 32'h1101b775;
         372:    rdata = 32'h4611cc22;
         373:    rdata = 32'h0048842a;
         374:    rdata = 32'h3f79ce06;
         375:    rdata = 32'h3d6d0048;
         376:    rdata = 32'h852285aa;
         377:    rdata = 32'h40f23f05;
         378:    rdata = 32'h61054462;
         379:    rdata = 32'h07938082;
         380:    rdata = 32'h06060300;
         381:    rdata = 32'h0ff67613;
         382:    rdata = 32'h00f50023;
         383:    rdata = 32'h07800793;
         384:    rdata = 32'h00f500a3;
         385:    rdata = 32'h87b24825;
         386:    rdata = 32'hf713c385;
         387:    rdata = 32'h069300f5;
         388:    rdata = 32'h64630577;
         389:    rdata = 32'h069300e8;
         390:    rdata = 32'h07330307;
         391:    rdata = 32'h00a300f5;
         392:    rdata = 32'h819100d7;
         393:    rdata = 32'hb7cd17fd;
         394:    rdata = 32'h01239532;
         395:    rdata = 32'h80820005;
         396:    rdata = 32'hbf754605;
         397:    rdata = 32'hbf654611;
         398:    rdata = 32'hcc221101;
         399:    rdata = 32'h842ace06;
         400:    rdata = 32'h0205d563;
         401:    rdata = 32'h02d00713;
         402:    rdata = 32'h00e50023;
         403:    rdata = 32'h40b005b3;
         404:    rdata = 32'h00484611;
         405:    rdata = 32'h00483715;
         406:    rdata = 32'h85aa3581;
         407:    rdata = 32'h00140513;
         408:    rdata = 32'h40f23d55;
         409:    rdata = 32'h61054462;
         410:    rdata = 32'h46118082;
         411:    rdata = 32'h37290048;
         412:    rdata = 32'h351d0048;
         413:    rdata = 32'h852285aa;
         414:    rdata = 32'h1141b7e5;
         415:    rdata = 32'hc606c422;
         416:    rdata = 32'h3535842a;
         417:    rdata = 32'h4703e115;
         418:    rdata = 32'h07930004;
         419:    rdata = 32'h1d630300;
         420:    rdata = 32'h470300f7;
         421:    rdata = 32'h07930014;
         422:    rdata = 32'h17630780;
         423:    rdata = 32'h852200f7;
         424:    rdata = 32'h40b24422;
         425:    rdata = 32'hbd250141;
         426:    rdata = 32'h442240b2;
         427:    rdata = 32'h80820141;
         428:    rdata = 32'hc4221141;
         429:    rdata = 32'h842ac606;
         430:    rdata = 32'h47833bdd;
         431:    rdata = 32'hc91d0004;
         432:    rdata = 32'h02d00693;
         433:    rdata = 32'h94634701;
         434:    rdata = 32'h872a00d7;
         435:    rdata = 32'h45010405;
         436:    rdata = 32'h46834629;
         437:    rdata = 32'hca810004;
         438:    rdata = 32'h02c507b3;
         439:    rdata = 32'hfd068513;
         440:    rdata = 32'h953e0405;
         441:    rdata = 32'hc319b7fd;
         442:    rdata = 32'h40a00533;
         443:    rdata = 32'h442240b2;
         444:    rdata = 32'h80820141;
         445:    rdata = 32'h03000713;
         446:    rdata = 32'h04e79663;
         447:    rdata = 32'h00144703;
         448:    rdata = 32'h07800793;
         449:    rdata = 32'h04f71063;
         450:    rdata = 32'h3bd18522;
         451:    rdata = 32'h0409cd05;
         452:    rdata = 32'h07134501;
         453:    rdata = 32'h06930600;
         454:    rdata = 32'h47830400;
         455:    rdata = 32'hd7f90004;
         456:    rdata = 32'h00f77a63;
         457:    rdata = 32'hfa978793;
         458:    rdata = 32'h0ff7f793;
         459:    rdata = 32'h8d5d0512;
         460:    rdata = 32'hb7e50405;
         461:    rdata = 32'h00f6f563;
         462:    rdata = 32'hfc978793;
         463:    rdata = 32'h8793b7f5;
         464:    rdata = 32'hb7ddfd07;
         465:    rdata = 32'hdeadc537;
         466:    rdata = 32'heef50513;
         467:    rdata = 32'h7793b745;
         468:    rdata = 32'h8793fdf5;
         469:    rdata = 32'hf793fbf7;
         470:    rdata = 32'h47650ff7;
         471:    rdata = 32'h00f77763;
         472:    rdata = 32'hfd050513;
         473:    rdata = 32'h00a53513;
         474:    rdata = 32'h45058082;
         475:    rdata = 32'hc10c8082;
         476:    rdata = 32'h8082c150;
         477:    rdata = 32'h99f14108;
         478:    rdata = 32'h8082952e;
         479:    rdata = 32'h80824148;
         480:    rdata = 32'hb0002573;
         481:    rdata = 32'hb80025f3;
         482:    rdata = 32'h00018082;
         483:    rdata = 32'h00010001;
         484:    rdata = 32'h00010001;
         485:    rdata = 32'h15fd0001;
         486:    rdata = 32'h8082f9ed;
         487:    rdata = 32'h8082c10c;
         488:    rdata = 32'h300462f3;
         489:    rdata = 32'h72f38082;
         490:    rdata = 32'h80823004;
         491:    rdata = 32'h62c1c14c;
         492:    rdata = 32'h3042a2f3;
         493:    rdata = 32'h22238082;
         494:    rdata = 32'h62c10005;
         495:    rdata = 32'h3042b2f3;
         496:    rdata = 32'hc50c8082;
         497:    rdata = 32'h000202b7;
         498:    rdata = 32'h3042a2f3;
         499:    rdata = 32'h24238082;
         500:    rdata = 32'h02b70005;
         501:    rdata = 32'hb2f30002;
         502:    rdata = 32'h80823042;
         503:    rdata = 32'hcc3e7139;
         504:    rdata = 32'hdc16de06;
         505:    rdata = 32'hd81eda1a;
         506:    rdata = 32'hd42ed62a;
         507:    rdata = 32'hd036d232;
         508:    rdata = 32'hca42ce3a;
         509:    rdata = 32'hc672c846;
         510:    rdata = 32'hc27ac476;
         511:    rdata = 32'h0797c07e;
         512:    rdata = 32'ha7830010;
         513:    rdata = 32'hc78d8027;
         514:    rdata = 32'h50f29782;
         515:    rdata = 32'h535252e2;
         516:    rdata = 32'h553253c2;
         517:    rdata = 32'h561255a2;
         518:    rdata = 32'h47725682;
         519:    rdata = 32'h485247e2;
         520:    rdata = 32'h4e3248c2;
         521:    rdata = 32'h4f124ea2;
         522:    rdata = 32'h61214f82;
         523:    rdata = 32'h30200073;
         524:    rdata = 32'h7139a001;
         525:    rdata = 32'hde06cc3e;
         526:    rdata = 32'hda1adc16;
         527:    rdata = 32'hd62ad81e;
         528:    rdata = 32'hd232d42e;
         529:    rdata = 32'hce3ad036;
         530:    rdata = 32'hc846ca42;
         531:    rdata = 32'hc476c672;
         532:    rdata = 32'hc07ec27a;
         533:    rdata = 32'h000ff797;
         534:    rdata = 32'h7b07a783;
         535:    rdata = 32'h50f29782;
         536:    rdata = 32'h535252e2;
         537:    rdata = 32'h553253c2;
         538:    rdata = 32'h561255a2;
         539:    rdata = 32'h47725682;
         540:    rdata = 32'h485247e2;
         541:    rdata = 32'h4e3248c2;
         542:    rdata = 32'h4f124ea2;
         543:    rdata = 32'h61214f82;
         544:    rdata = 32'h30200073;
         545:    rdata = 32'hcc3e7139;
         546:    rdata = 32'hdc16de06;
         547:    rdata = 32'hd81eda1a;
         548:    rdata = 32'hd42ed62a;
         549:    rdata = 32'hd036d232;
         550:    rdata = 32'hca42ce3a;
         551:    rdata = 32'hc672c846;
         552:    rdata = 32'hc27ac476;
         553:    rdata = 32'hf797c07e;
         554:    rdata = 32'ha783000f;
         555:    rdata = 32'h97827627;
         556:    rdata = 32'h52e250f2;
         557:    rdata = 32'h53c25352;
         558:    rdata = 32'h55a25532;
         559:    rdata = 32'h56825612;
         560:    rdata = 32'h47e24772;
         561:    rdata = 32'h48c24852;
         562:    rdata = 32'h4ea24e32;
         563:    rdata = 32'h4f824f12;
         564:    rdata = 32'h00736121;
         565:    rdata = 32'h87933020;
         566:    rdata = 32'hc15c0045;
         567:    rdata = 32'h00858793;
         568:    rdata = 32'h8793c51c;
         569:    rdata = 32'hc55c00c5;
         570:    rdata = 32'h01058793;
         571:    rdata = 32'h8793c91c;
         572:    rdata = 32'hc95c0145;
         573:    rdata = 32'h01858793;
         574:    rdata = 32'hcd1cc10c;
         575:    rdata = 32'h01c58793;
         576:    rdata = 32'h02058593;
         577:    rdata = 32'hd10ccd5c;
         578:    rdata = 32'h511c8082;
         579:    rdata = 32'h16338a05;
         580:    rdata = 32'h439c00b6;
         581:    rdata = 32'h48b797b3;
         582:    rdata = 32'h511c8e5d;
         583:    rdata = 32'h8082c390;
         584:    rdata = 32'h4388511c;
         585:    rdata = 32'h97b34785;
         586:    rdata = 32'h8d7d00b7;
         587:    rdata = 32'h00a03533;
         588:    rdata = 32'h455c8082;
         589:    rdata = 32'h47854388;
         590:    rdata = 32'h00b797b3;
         591:    rdata = 32'h35338d7d;
         592:    rdata = 32'h808200a0;
         593:    rdata = 32'h439c451c;
         594:    rdata = 32'h8e6d8e3d;
         595:    rdata = 32'h451c8e3d;
         596:    rdata = 32'h8082c390;
         597:    rdata = 32'h16334785;
         598:    rdata = 32'h95b300b6;
         599:    rdata = 32'hb7dd00b7;
         600:    rdata = 32'hc4221141;
         601:    rdata = 32'hc606c226;
         602:    rdata = 32'h84ae842a;
         603:    rdata = 32'h461337d9;
         604:    rdata = 32'h85220015;
         605:    rdata = 32'h40b24422;
         606:    rdata = 32'h449285a6;
         607:    rdata = 32'h0ff67613;
         608:    rdata = 32'hbfc90141;
         609:    rdata = 32'h4388455c;
         610:    rdata = 32'h49155513;
         611:    rdata = 32'h455c8082;
         612:    rdata = 32'h55134388;
         613:    rdata = 32'h80824905;
         614:    rdata = 32'hc2261141;
         615:    rdata = 32'h84ae4601;
         616:    rdata = 32'hc42245bd;
         617:    rdata = 32'h842ac606;
         618:    rdata = 32'h8522378d;
         619:    rdata = 32'h40b24422;
         620:    rdata = 32'h44928626;
         621:    rdata = 32'h014145bd;
         622:    rdata = 32'h8793bf71;
         623:    rdata = 32'hc15c0045;
         624:    rdata = 32'h00858793;
         625:    rdata = 32'hc51cc10c;
         626:    rdata = 32'h00c58793;
         627:    rdata = 32'hc55c05c1;
         628:    rdata = 32'h8082c90c;
         629:    rdata = 32'hf7934118;
         630:    rdata = 32'h430c0015;
         631:    rdata = 32'h8ddd99f9;
         632:    rdata = 32'h8082c30c;
         633:    rdata = 32'h89854118;
         634:    rdata = 32'h00159793;
         635:    rdata = 32'h99f5430c;
         636:    rdata = 32'hc30c8ddd;
         637:    rdata = 32'h491c8082;
         638:    rdata = 32'h00b78023;
         639:    rdata = 32'h451c8082;
         640:    rdata = 32'h00078023;
         641:    rdata = 32'h439c415c;
         642:    rdata = 32'hdfed8b85;
         643:    rdata = 32'hc503455c;
         644:    rdata = 32'h75130007;
         645:    rdata = 32'h80820ff5;
         646:    rdata = 32'h8023451c;
         647:    rdata = 32'h415c00b7;
         648:    rdata = 32'hd793439c;
         649:    rdata = 32'hffe54817;
         650:    rdata = 32'hc783455c;
         651:    rdata = 32'h80820007;
         652:    rdata = 32'h4388415c;
         653:    rdata = 32'h80828905;
         654:    rdata = 32'h4388415c;
         655:    rdata = 32'h48155513;
         656:    rdata = 32'h87938082;
         657:    rdata = 32'hc15c0045;
         658:    rdata = 32'h00858793;
         659:    rdata = 32'h8793c51c;
         660:    rdata = 32'hc55c00c5;
         661:    rdata = 32'h01058793;
         662:    rdata = 32'h47b1c91c;
         663:    rdata = 32'h8823c10c;
         664:    rdata = 32'h419c00f5;
         665:    rdata = 32'h0017e793;
         666:    rdata = 32'h8082c19c;
         667:    rdata = 32'h439c415c;
         668:    rdata = 32'hdfed8b85;
         669:    rdata = 32'hc503455c;
         670:    rdata = 32'h75130007;
         671:    rdata = 32'h80820ff5;
         672:    rdata = 32'hcc221101;
         673:    rdata = 32'hc84aca26;
         674:    rdata = 32'hc256c64e;
         675:    rdata = 32'hce06c05a;
         676:    rdata = 32'h84aac452;
         677:    rdata = 32'h89b2892e;
         678:    rdata = 32'h4aa94401;
         679:    rdata = 32'h5f634b21;
         680:    rdata = 32'h85260334;
         681:    rdata = 32'h00890a33;
         682:    rdata = 32'h002337d1;
         683:    rdata = 32'h1f6300aa;
         684:    rdata = 32'h00230155;
         685:    rdata = 32'h4501000a;
         686:    rdata = 32'h446240f2;
         687:    rdata = 32'h494244d2;
         688:    rdata = 32'h4a2249b2;
         689:    rdata = 32'h4b024a92;
         690:    rdata = 32'h80826105;
         691:    rdata = 32'h01651463;
         692:    rdata = 32'h1479c401;
         693:    rdata = 32'hb7e10405;
         694:    rdata = 32'hbfed547d;
         695:    rdata = 32'hbfe94505;
         696:    rdata = 32'h8023451c;
         697:    rdata = 32'h415c00b7;
         698:    rdata = 32'hd793439c;
         699:    rdata = 32'hffe54817;
         700:    rdata = 32'h11418082;
         701:    rdata = 32'hc226c422;
         702:    rdata = 32'h84aac606;
         703:    rdata = 32'h4583842e;
         704:    rdata = 32'hc5890004;
         705:    rdata = 32'h04058526;
         706:    rdata = 32'hbfd53fe1;
         707:    rdata = 32'h442240b2;
         708:    rdata = 32'h01414492;
         709:    rdata = 32'h415c8082;
         710:    rdata = 32'h89054388;
         711:    rdata = 32'h455c8082;
         712:    rdata = 32'h0007c503;
         713:    rdata = 32'h0ff57513;
         714:    rdata = 32'h11418082;
         715:    rdata = 32'h00000597;
         716:    rdata = 32'h14c58593;
         717:    rdata = 32'h000ff517;
         718:    rdata = 32'h52450513;
         719:    rdata = 32'hf0efc606;
         720:    rdata = 32'hf0ef8bdf;
         721:    rdata = 32'hf517f82f;
         722:    rdata = 32'h0513000f;
         723:    rdata = 32'h3d1d4c65;
         724:    rdata = 32'h0597c121;
         725:    rdata = 32'h85930000;
         726:    rdata = 32'hf5171425;
         727:    rdata = 32'h0513000f;
         728:    rdata = 32'hf0ef4fe5;
         729:    rdata = 32'h62c1899f;
         730:    rdata = 32'h305292f3;
         731:    rdata = 32'h00000597;
         732:    rdata = 32'h1bc58593;
         733:    rdata = 32'h000ff517;
         734:    rdata = 32'h4e450513;
         735:    rdata = 32'h87fff0ef;
         736:    rdata = 32'h801ff0ef;
         737:    rdata = 32'h4fc0f06f;
         738:    rdata = 32'h450140b2;
         739:    rdata = 32'h80820141;
         740:    rdata = 32'h000ff517;
         741:    rdata = 32'h47c50513;
         742:    rdata = 32'hc5393bdd;
         743:    rdata = 32'h00000597;
         744:    rdata = 32'h11058593;
         745:    rdata = 32'h000ff517;
         746:    rdata = 32'h4b450513;
         747:    rdata = 32'h84fff0ef;
         748:    rdata = 32'he5eff0ef;
         749:    rdata = 32'h0597cd09;
         750:    rdata = 32'h85930000;
         751:    rdata = 32'hf5171165;
         752:    rdata = 32'h0513000f;
         753:    rdata = 32'hf0ef49a5;
         754:    rdata = 32'hf0ef835f;
         755:    rdata = 32'h0597f88f;
         756:    rdata = 32'h85930000;
         757:    rdata = 32'hf51713e5;
         758:    rdata = 32'h0513000f;
         759:    rdata = 32'hf0ef4825;
         760:    rdata = 32'hf0ef81df;
         761:    rdata = 32'hb741f14f;
         762:    rdata = 32'h00000597;
         763:    rdata = 32'h10858593;
         764:    rdata = 32'h000ff517;
         765:    rdata = 32'h46850513;
         766:    rdata = 32'h803ff0ef;
         767:    rdata = 32'hd98ff0ef;
         768:    rdata = 32'hf797b7f9;
         769:    rdata = 32'h8793000f;
         770:    rdata = 32'h674145a7;
         771:    rdata = 32'h6711c398;
         772:    rdata = 32'h8082c3d8;
         773:    rdata = 32'h010005b7;
         774:    rdata = 32'h000ff517;
         775:    rdata = 32'h3f450513;
         776:    rdata = 32'h17b7b95d;
         777:    rdata = 32'hf7170100;
         778:    rdata = 32'h0713000f;
         779:    rdata = 32'h869340a7;
         780:    rdata = 32'hc3540047;
         781:    rdata = 32'h00878693;
         782:    rdata = 32'hc714c31c;
         783:    rdata = 32'h00c78693;
         784:    rdata = 32'hc75407c1;
         785:    rdata = 32'h8082cb1c;
         786:    rdata = 32'h010025b7;
         787:    rdata = 32'h000ff517;
         788:    rdata = 32'h3f850513;
         789:    rdata = 32'h0000b3fd;
         790:    rdata = 32'h00000000;
         791:    rdata = 32'h00000000;
         792:    rdata = 32'h00000000;
         793:    rdata = 32'h00000000;
         794:    rdata = 32'h00000c02;
         795:    rdata = 32'h00000c14;
         796:    rdata = 32'h00000c22;
         797:    rdata = 32'h00000c48;
         798:    rdata = 32'h4f464e49;
         799:    rdata = 32'h6f62203a;
         800:    rdata = 32'h6f6c746f;
         801:    rdata = 32'h72656461;
         802:    rdata = 32'h61747320;
         803:    rdata = 32'h64657472;
         804:    rdata = 32'h0000000a;
         805:    rdata = 32'h4f464e49;
         806:    rdata = 32'h6f63203a;
         807:    rdata = 32'h6f6c6564;
         808:    rdata = 32'h73206461;
         809:    rdata = 32'h7070696b;
         810:    rdata = 32'h000a6465;
         811:    rdata = 32'h4f464e49;
         812:    rdata = 32'h6f63203a;
         813:    rdata = 32'h6f6c6564;
         814:    rdata = 32'h73206461;
         815:    rdata = 32'h6372756f;
         816:    rdata = 32'h75203a65;
         817:    rdata = 32'h0a747261;
         818:    rdata = 32'h00000000;
         819:    rdata = 32'h4f525245;
         820:    rdata = 32'h63203a52;
         821:    rdata = 32'h6c65646f;
         822:    rdata = 32'h2064616f;
         823:    rdata = 32'h656d6974;
         824:    rdata = 32'h2074756f;
         825:    rdata = 32'h7563636f;
         826:    rdata = 32'h64657272;
         827:    rdata = 32'h0000000a;
         828:    rdata = 32'h4f464e49;
         829:    rdata = 32'h6f63203a;
         830:    rdata = 32'h6f6c6564;
         831:    rdata = 32'h73206461;
         832:    rdata = 32'h6372756f;
         833:    rdata = 32'h73203a65;
         834:    rdata = 32'h000a6970;
         835:    rdata = 32'h4f464e49;
         836:    rdata = 32'h6f63203a;
         837:    rdata = 32'h6f6c6564;
         838:    rdata = 32'h66206461;
         839:    rdata = 32'h73696e69;
         840:    rdata = 32'h0a646568;
         841:    rdata = 32'h00000000;
         842:    rdata = 32'h4f464e49;
         843:    rdata = 32'h6f62203a;
         844:    rdata = 32'h6f6c746f;
         845:    rdata = 32'h72656461;
         846:    rdata = 32'h6e696620;
         847:    rdata = 32'h65687369;
         848:    rdata = 32'h00000a64;
         849:    rdata = 32'h0000203a;
         850:    rdata = 32'h6f636e69;
         851:    rdata = 32'h63657272;
         852:    rdata = 32'h61762074;
         853:    rdata = 32'h2e65756c;
         854:    rdata = 32'h79727420;
         855:    rdata = 32'h61676120;
         856:    rdata = 32'h000a6e69;
        default: rdata = 32'h00000000;
    endcase
end
endmodule
