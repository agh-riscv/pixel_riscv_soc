/**
 * Copyright (C) 2020  AGH University of Science and Technology
 *
 * This program is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with this program.  If not, see <https://www.gnu.org/licenses/>.
 */

module spi_mem (
    output logic [31:0] rdata,
    input logic [31:0] addr
);

/**
 * Module internal logic
 */

always_comb begin
    case (addr[13:2])
           0:    rdata = 32'h15e0006f;
           1:    rdata = 32'h15a0006f;
           2:    rdata = 32'h1560006f;
           3:    rdata = 32'h1520006f;
           4:    rdata = 32'h14e0006f;
           5:    rdata = 32'h14a0006f;
           6:    rdata = 32'h1460006f;
           7:    rdata = 32'h1420006f;
           8:    rdata = 32'h13e0006f;
           9:    rdata = 32'h13a0006f;
          10:    rdata = 32'h1360006f;
          11:    rdata = 32'h1320006f;
          12:    rdata = 32'h12e0006f;
          13:    rdata = 32'h12a0006f;
          14:    rdata = 32'h1260006f;
          15:    rdata = 32'h1220006f;
          16:    rdata = 32'h04c0006f;
          17:    rdata = 32'h0a80006f;
          18:    rdata = 32'h1160006f;
          19:    rdata = 32'h1120006f;
          20:    rdata = 32'h10e0006f;
          21:    rdata = 32'h10a0006f;
          22:    rdata = 32'h1060006f;
          23:    rdata = 32'h1020006f;
          24:    rdata = 32'h0fe0006f;
          25:    rdata = 32'h0fa0006f;
          26:    rdata = 32'h0f60006f;
          27:    rdata = 32'h0f20006f;
          28:    rdata = 32'h0ee0006f;
          29:    rdata = 32'h0ea0006f;
          30:    rdata = 32'h0e60006f;
          31:    rdata = 32'h0e20006f;
          32:    rdata = 32'h0e20006f;
          33:    rdata = 32'h0da0006f;
          34:    rdata = 32'h0d60006f;
          35:    rdata = 32'hde22715d;
          36:    rdata = 32'h01000437;
          37:    rdata = 32'h484cda2e;
          38:    rdata = 32'h0517dc2a;
          39:    rdata = 32'h05130000;
          40:    rdata = 32'hc6864fa5;
          41:    rdata = 32'hc29ac496;
          42:    rdata = 32'hd832c09e;
          43:    rdata = 32'hd43ad636;
          44:    rdata = 32'hd042d23e;
          45:    rdata = 32'hcc72ce46;
          46:    rdata = 32'hc87aca76;
          47:    rdata = 32'h2611c67e;
          48:    rdata = 32'h00042a23;
          49:    rdata = 32'h40b65472;
          50:    rdata = 32'h431642a6;
          51:    rdata = 32'h55624386;
          52:    rdata = 32'h564255d2;
          53:    rdata = 32'h572256b2;
          54:    rdata = 32'h58025792;
          55:    rdata = 32'h4e6248f2;
          56:    rdata = 32'h4f424ed2;
          57:    rdata = 32'h61614fb2;
          58:    rdata = 32'h30200073;
          59:    rdata = 32'hde22715d;
          60:    rdata = 32'h000f0417;
          61:    rdata = 32'hf1040413;
          62:    rdata = 32'h4583da2e;
          63:    rdata = 32'hdc2a0004;
          64:    rdata = 32'hd43a4505;
          65:    rdata = 32'hc686d23e;
          66:    rdata = 32'hc29ac496;
          67:    rdata = 32'hd832c09e;
          68:    rdata = 32'hd042d636;
          69:    rdata = 32'hcc72ce46;
          70:    rdata = 32'hc87aca76;
          71:    rdata = 32'h2215c67e;
          72:    rdata = 32'h00044783;
          73:    rdata = 32'h01003737;
          74:    rdata = 32'h0017c793;
          75:    rdata = 32'h00f40023;
          76:    rdata = 32'h9bf9435c;
          77:    rdata = 32'h5472c35c;
          78:    rdata = 32'h42a640b6;
          79:    rdata = 32'h43864316;
          80:    rdata = 32'h55d25562;
          81:    rdata = 32'h56b25642;
          82:    rdata = 32'h57925722;
          83:    rdata = 32'h48f25802;
          84:    rdata = 32'h4ed24e62;
          85:    rdata = 32'h4fb24f42;
          86:    rdata = 32'h00736161;
          87:    rdata = 32'h006f3020;
          88:    rdata = 32'h00930000;
          89:    rdata = 32'h01130000;
          90:    rdata = 32'h01930000;
          91:    rdata = 32'h02130000;
          92:    rdata = 32'h02930000;
          93:    rdata = 32'h03130000;
          94:    rdata = 32'h03930000;
          95:    rdata = 32'h04130000;
          96:    rdata = 32'h04930000;
          97:    rdata = 32'h05130000;
          98:    rdata = 32'h05930000;
          99:    rdata = 32'h06130000;
         100:    rdata = 32'h06930000;
         101:    rdata = 32'h07130000;
         102:    rdata = 32'h07930000;
         103:    rdata = 32'h08130000;
         104:    rdata = 32'h08930000;
         105:    rdata = 32'h09130000;
         106:    rdata = 32'h09930000;
         107:    rdata = 32'h0a130000;
         108:    rdata = 32'h0a930000;
         109:    rdata = 32'h0b130000;
         110:    rdata = 32'h0b930000;
         111:    rdata = 32'h0c130000;
         112:    rdata = 32'h0c930000;
         113:    rdata = 32'h0d130000;
         114:    rdata = 32'h0d930000;
         115:    rdata = 32'h0e130000;
         116:    rdata = 32'h0e930000;
         117:    rdata = 32'h0f130000;
         118:    rdata = 32'h0f930000;
         119:    rdata = 32'h41170000;
         120:    rdata = 32'h0113000f;
         121:    rdata = 32'h0297e221;
         122:    rdata = 32'h8293000f;
         123:    rdata = 32'h0317e1a2;
         124:    rdata = 32'h0313000f;
         125:    rdata = 32'hd863e133;
         126:    rdata = 32'ha0230062;
         127:    rdata = 32'h82930002;
         128:    rdata = 32'h5ce30042;
         129:    rdata = 32'h0297fe53;
         130:    rdata = 32'h82930000;
         131:    rdata = 32'h03173ba2;
         132:    rdata = 32'h0313000f;
         133:    rdata = 32'h0397df23;
         134:    rdata = 32'h8393000f;
         135:    rdata = 32'h5c63dea3;
         136:    rdata = 32'hae030073;
         137:    rdata = 32'h20230002;
         138:    rdata = 32'h829301c3;
         139:    rdata = 32'h03130042;
         140:    rdata = 32'hd8e30043;
         141:    rdata = 32'h0513fe63;
         142:    rdata = 32'h05930000;
         143:    rdata = 32'h00ef0000;
         144:    rdata = 32'h07b73000;
         145:    rdata = 32'h47980100;
         146:    rdata = 32'h8de98db9;
         147:    rdata = 32'hc78c8db9;
         148:    rdata = 32'h62f38082;
         149:    rdata = 32'h80823004;
         150:    rdata = 32'ha2f362c1;
         151:    rdata = 32'h80823042;
         152:    rdata = 32'h000202b7;
         153:    rdata = 32'h3042a2f3;
         154:    rdata = 32'h80828082;
         155:    rdata = 32'h27b78082;
         156:    rdata = 32'h47190100;
         157:    rdata = 32'h00e78823;
         158:    rdata = 32'h67134398;
         159:    rdata = 32'hc3980017;
         160:    rdata = 32'h27378082;
         161:    rdata = 32'h435c0100;
         162:    rdata = 32'hdff58b85;
         163:    rdata = 32'h00c74503;
         164:    rdata = 32'h0ff57513;
         165:    rdata = 32'h11018082;
         166:    rdata = 32'hca26cc22;
         167:    rdata = 32'hc452c84a;
         168:    rdata = 32'hc64ece06;
         169:    rdata = 32'h84ae892a;
         170:    rdata = 32'h4a294401;
         171:    rdata = 32'h00944463;
         172:    rdata = 32'ha8194505;
         173:    rdata = 32'h008909b3;
         174:    rdata = 32'h802337e9;
         175:    rdata = 32'h1d6300a9;
         176:    rdata = 32'h80230145;
         177:    rdata = 32'h45010009;
         178:    rdata = 32'h446240f2;
         179:    rdata = 32'h494244d2;
         180:    rdata = 32'h4a2249b2;
         181:    rdata = 32'h80826105;
         182:    rdata = 32'hbfc90405;
         183:    rdata = 32'h010027b7;
         184:    rdata = 32'h00a78423;
         185:    rdata = 32'h01002737;
         186:    rdata = 32'hd793435c;
         187:    rdata = 32'hffed4817;
         188:    rdata = 32'h11418082;
         189:    rdata = 32'hc606c422;
         190:    rdata = 32'h4503842a;
         191:    rdata = 32'he5110004;
         192:    rdata = 32'h40b24422;
         193:    rdata = 32'h01414529;
         194:    rdata = 32'h0405bfd1;
         195:    rdata = 32'hb7f53fc1;
         196:    rdata = 32'hdca27119;
         197:    rdata = 32'h85aa842e;
         198:    rdata = 32'hde860068;
         199:    rdata = 32'h0597228d;
         200:    rdata = 32'h85930000;
         201:    rdata = 32'h00682965;
         202:    rdata = 32'h85a222a5;
         203:    rdata = 32'h228d0068;
         204:    rdata = 32'h37c10068;
         205:    rdata = 32'h546650f6;
         206:    rdata = 32'h80826109;
         207:    rdata = 32'hdaa67119;
         208:    rdata = 32'h85aa84ae;
         209:    rdata = 32'hde860068;
         210:    rdata = 32'h8432dca2;
         211:    rdata = 32'h05972a0d;
         212:    rdata = 32'h85930000;
         213:    rdata = 32'h006826a5;
         214:    rdata = 32'h85a62a25;
         215:    rdata = 32'h2a0d0068;
         216:    rdata = 32'h00000597;
         217:    rdata = 32'h25c58593;
         218:    rdata = 32'h221d0068;
         219:    rdata = 32'h006885a2;
         220:    rdata = 32'h00682205;
         221:    rdata = 32'h50f63fbd;
         222:    rdata = 32'h54d65466;
         223:    rdata = 32'h80826109;
         224:    rdata = 32'h85aa1101;
         225:    rdata = 32'hce060048;
         226:    rdata = 32'h00482ab1;
         227:    rdata = 32'h40f2379d;
         228:    rdata = 32'h80826105;
         229:    rdata = 32'h85aa1101;
         230:    rdata = 32'hce060048;
         231:    rdata = 32'h00482a11;
         232:    rdata = 32'h40f23f89;
         233:    rdata = 32'h80826105;
         234:    rdata = 32'hcc221101;
         235:    rdata = 32'h0048842a;
         236:    rdata = 32'h2a0dce06;
         237:    rdata = 32'h8522004c;
         238:    rdata = 32'h40f23fa1;
         239:    rdata = 32'h61054462;
         240:    rdata = 32'h11018082;
         241:    rdata = 32'h842acc22;
         242:    rdata = 32'hce060048;
         243:    rdata = 32'h004c20d5;
         244:    rdata = 32'h3f3d8522;
         245:    rdata = 32'h446240f2;
         246:    rdata = 32'h80826105;
         247:    rdata = 32'hd4227179;
         248:    rdata = 32'h0028842a;
         249:    rdata = 32'hd226d606;
         250:    rdata = 32'h20d984b2;
         251:    rdata = 32'h084885a6;
         252:    rdata = 32'h085028d5;
         253:    rdata = 32'h8522002c;
         254:    rdata = 32'h50b23791;
         255:    rdata = 32'h54925422;
         256:    rdata = 32'h80826145;
         257:    rdata = 32'hd4227179;
         258:    rdata = 32'h0028842a;
         259:    rdata = 32'hd226d606;
         260:    rdata = 32'h287984b2;
         261:    rdata = 32'h084885a6;
         262:    rdata = 32'h08502861;
         263:    rdata = 32'h8522002c;
         264:    rdata = 32'h50b23f31;
         265:    rdata = 32'h54925422;
         266:    rdata = 32'h80826145;
         267:    rdata = 32'h03000793;
         268:    rdata = 32'h76130606;
         269:    rdata = 32'h00230ff6;
         270:    rdata = 32'h079300f5;
         271:    rdata = 32'h00a30780;
         272:    rdata = 32'h079300f5;
         273:    rdata = 32'hf7930016;
         274:    rdata = 32'h97aa0ff7;
         275:    rdata = 32'h00150693;
         276:    rdata = 32'hf7134825;
         277:    rdata = 32'h616300f5;
         278:    rdata = 32'h071302e8;
         279:    rdata = 32'h80230307;
         280:    rdata = 32'h17fd00e7;
         281:    rdata = 32'h96e38191;
         282:    rdata = 32'h0609fef6;
         283:    rdata = 32'h0ff67613;
         284:    rdata = 32'h0023962a;
         285:    rdata = 32'h80820006;
         286:    rdata = 32'h05770713;
         287:    rdata = 32'h87aab7cd;
         288:    rdata = 32'h0005c703;
         289:    rdata = 32'h07850585;
         290:    rdata = 32'hfee78fa3;
         291:    rdata = 32'h8082fb75;
         292:    rdata = 32'hc68387aa;
         293:    rdata = 32'h873e0007;
         294:    rdata = 32'hfee50785;
         295:    rdata = 32'h0005c783;
         296:    rdata = 32'h07050585;
         297:    rdata = 32'hfef70fa3;
         298:    rdata = 32'h8082fbf5;
         299:    rdata = 32'hbfbd4605;
         300:    rdata = 32'hbfad4611;
         301:    rdata = 32'h00350613;
         302:    rdata = 32'h06400793;
         303:    rdata = 32'hd7334829;
         304:    rdata = 32'h050502f5;
         305:    rdata = 32'h0ff77693;
         306:    rdata = 32'h02f686b3;
         307:    rdata = 32'h03070713;
         308:    rdata = 32'hfee50fa3;
         309:    rdata = 32'h0307d7b3;
         310:    rdata = 32'h12e38d95;
         311:    rdata = 32'h0023fea6;
         312:    rdata = 32'h80820006;
         313:    rdata = 32'h00581101;
         314:    rdata = 32'h3b9ad7b7;
         315:    rdata = 32'hce0686ae;
         316:    rdata = 32'ha0078793;
         317:    rdata = 32'h432985ba;
         318:    rdata = 32'h00e10893;
         319:    rdata = 32'h02f6d633;
         320:    rdata = 32'h78130705;
         321:    rdata = 32'h08330ff6;
         322:    rdata = 32'h061302f8;
         323:    rdata = 32'h0fa30306;
         324:    rdata = 32'hd7b3fec7;
         325:    rdata = 32'h86b30267;
         326:    rdata = 32'h11e34106;
         327:    rdata = 32'h0723ff17;
         328:    rdata = 32'h07130001;
         329:    rdata = 32'hc7830300;
         330:    rdata = 32'h88630005;
         331:    rdata = 32'he39100e7;
         332:    rdata = 32'h37b115fd;
         333:    rdata = 32'h610540f2;
         334:    rdata = 32'h05858082;
         335:    rdata = 32'h7119b7ed;
         336:    rdata = 32'h3335de86;
         337:    rdata = 32'h00000517;
         338:    rdata = 32'h05c50513;
         339:    rdata = 32'h07b7335d;
         340:    rdata = 32'h473d0100;
         341:    rdata = 32'hcf98cb98;
         342:    rdata = 32'h33193301;
         343:    rdata = 32'hf73739dd;
         344:    rdata = 32'h37b702fa;
         345:    rdata = 32'h07130100;
         346:    rdata = 32'hc7d807f7;
         347:    rdata = 32'h67134398;
         348:    rdata = 32'hc3980017;
         349:    rdata = 32'h06400593;
         350:    rdata = 32'h3b310068;
         351:    rdata = 32'h3b950068;
         352:    rdata = 32'h0000bfd5;
         353:    rdata = 32'h00000000;
         354:    rdata = 32'h00000000;
         355:    rdata = 32'h00000000;
         356:    rdata = 32'h00000000;
         357:    rdata = 32'h4f495047;
         358:    rdata = 32'h53493e2d;
         359:    rdata = 32'h00000052;
         360:    rdata = 32'h6c707061;
         361:    rdata = 32'h74616369;
         362:    rdata = 32'h206e6f69;
         363:    rdata = 32'h72617473;
         364:    rdata = 32'h00646574;
         365:    rdata = 32'h0000203a;
         366:    rdata = 32'h00002820;
         367:    rdata = 32'h00203a29;
        default: rdata = 32'h00000000;
    endcase
end
endmodule
