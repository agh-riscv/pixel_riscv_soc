/**
 * Copyright (C) 2020  AGH University of Science and Technology
 *
 * This program is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with this program.  If not, see <https://www.gnu.org/licenses/>.
 */

module spi_mem (
    output logic [31:0] rdata,
    input logic [31:0] addr
);

/**
 * Module internal logic
 */

always_comb begin
    case (addr[13:2])
           0:    rdata = 32'h24a0106f;
           1:    rdata = 32'h0880006f;
           2:    rdata = 32'h0840006f;
           3:    rdata = 32'h0800006f;
           4:    rdata = 32'h07c0006f;
           5:    rdata = 32'h0780006f;
           6:    rdata = 32'h0740006f;
           7:    rdata = 32'h0700006f;
           8:    rdata = 32'h06c0006f;
           9:    rdata = 32'h0680006f;
          10:    rdata = 32'h0640006f;
          11:    rdata = 32'h0600006f;
          12:    rdata = 32'h05c0006f;
          13:    rdata = 32'h0580006f;
          14:    rdata = 32'h0540006f;
          15:    rdata = 32'h0500006f;
          16:    rdata = 32'h2600106f;
          17:    rdata = 32'h2ae0106f;
          18:    rdata = 32'h0440006f;
          19:    rdata = 32'h0400006f;
          20:    rdata = 32'h03c0006f;
          21:    rdata = 32'h0380006f;
          22:    rdata = 32'h0340006f;
          23:    rdata = 32'h0300006f;
          24:    rdata = 32'h02c0006f;
          25:    rdata = 32'h0280006f;
          26:    rdata = 32'h0240006f;
          27:    rdata = 32'h0200006f;
          28:    rdata = 32'h01c0006f;
          29:    rdata = 32'h0180006f;
          30:    rdata = 32'h0140006f;
          31:    rdata = 32'h0100006f;
          32:    rdata = 32'h0100006f;
          33:    rdata = 32'h0080006f;
          34:    rdata = 32'h0040006f;
          35:    rdata = 32'h0000006f;
          36:    rdata = 32'h00000093;
          37:    rdata = 32'h00000113;
          38:    rdata = 32'h00000193;
          39:    rdata = 32'h00000213;
          40:    rdata = 32'h00000293;
          41:    rdata = 32'h00000313;
          42:    rdata = 32'h00000393;
          43:    rdata = 32'h00000413;
          44:    rdata = 32'h00000493;
          45:    rdata = 32'h00000513;
          46:    rdata = 32'h00000593;
          47:    rdata = 32'h00000613;
          48:    rdata = 32'h00000693;
          49:    rdata = 32'h00000713;
          50:    rdata = 32'h00000793;
          51:    rdata = 32'h00000813;
          52:    rdata = 32'h00000893;
          53:    rdata = 32'h00000913;
          54:    rdata = 32'h00000993;
          55:    rdata = 32'h00000a13;
          56:    rdata = 32'h00000a93;
          57:    rdata = 32'h00000b13;
          58:    rdata = 32'h00000b93;
          59:    rdata = 32'h00000c13;
          60:    rdata = 32'h00000c93;
          61:    rdata = 32'h00000d13;
          62:    rdata = 32'h00000d93;
          63:    rdata = 32'h00000e13;
          64:    rdata = 32'h00000e93;
          65:    rdata = 32'h00000f13;
          66:    rdata = 32'h00000f93;
          67:    rdata = 32'h000f4117;
          68:    rdata = 32'hef410113;
          69:    rdata = 32'h000f0297;
          70:    rdata = 32'heec28293;
          71:    rdata = 32'h000f0317;
          72:    rdata = 32'hf7830313;
          73:    rdata = 32'h0062d863;
          74:    rdata = 32'h0002a023;
          75:    rdata = 32'h00428293;
          76:    rdata = 32'hfe535ce3;
          77:    rdata = 32'h00002297;
          78:    rdata = 32'heb028293;
          79:    rdata = 32'h000f0317;
          80:    rdata = 32'hec430313;
          81:    rdata = 32'h000f0397;
          82:    rdata = 32'hebc38393;
          83:    rdata = 32'h00735c63;
          84:    rdata = 32'h0002ae03;
          85:    rdata = 32'h01c32023;
          86:    rdata = 32'h00428293;
          87:    rdata = 32'h00430313;
          88:    rdata = 32'hfe7348e3;
          89:    rdata = 32'h00002297;
          90:    rdata = 32'h86428293;
          91:    rdata = 32'h00002317;
          92:    rdata = 32'h87030313;
          93:    rdata = 32'h0062da63;
          94:    rdata = 32'h0002a783;
          95:    rdata = 32'h000780e7;
          96:    rdata = 32'h00428293;
          97:    rdata = 32'hfe62cae3;
          98:    rdata = 32'h00000513;
          99:    rdata = 32'h00000593;
         100:    rdata = 32'h7a0010ef;
         101:    rdata = 32'h25971141;
         102:    rdata = 32'h85930000;
         103:    rdata = 32'h051795e5;
         104:    rdata = 32'h0513000f;
         105:    rdata = 32'hc606eea5;
         106:    rdata = 32'h7a9000ef;
         107:    rdata = 32'h051740b2;
         108:    rdata = 32'h0513000f;
         109:    rdata = 32'h0141eb25;
         110:    rdata = 32'h47a0106f;
         111:    rdata = 32'h00002597;
         112:    rdata = 32'h94458593;
         113:    rdata = 32'h000f0517;
         114:    rdata = 32'hec450513;
         115:    rdata = 32'h7850006f;
         116:    rdata = 32'h00002597;
         117:    rdata = 32'hb8458593;
         118:    rdata = 32'h000f0517;
         119:    rdata = 32'heb050513;
         120:    rdata = 32'h7710006f;
         121:    rdata = 32'h00002597;
         122:    rdata = 32'hb9058593;
         123:    rdata = 32'h000f0517;
         124:    rdata = 32'he9c50513;
         125:    rdata = 32'h75d0006f;
         126:    rdata = 32'h114141d8;
         127:    rdata = 32'hc422c606;
         128:    rdata = 32'hc04ac226;
         129:    rdata = 32'hc4634785;
         130:    rdata = 32'h259702e7;
         131:    rdata = 32'h85930000;
         132:    rdata = 32'h0517b725;
         133:    rdata = 32'h0513000f;
         134:    rdata = 32'h00efe765;
         135:    rdata = 32'h44057370;
         136:    rdata = 32'h852240b2;
         137:    rdata = 32'h44924422;
         138:    rdata = 32'h01414902;
         139:    rdata = 32'h45808082;
         140:    rdata = 32'h146384ae;
         141:    rdata = 32'h519c00f4;
         142:    rdata = 32'h2597c791;
         143:    rdata = 32'h85930000;
         144:    rdata = 32'hbfc1b5e5;
         145:    rdata = 32'h02458913;
         146:    rdata = 32'h2597854a;
         147:    rdata = 32'h85930000;
         148:    rdata = 32'h00efb725;
         149:    rdata = 32'hc50d4970;
         150:    rdata = 32'h00002597;
         151:    rdata = 32'hb6858593;
         152:    rdata = 32'h00ef854a;
         153:    rdata = 32'hcd014870;
         154:    rdata = 32'h00002597;
         155:    rdata = 32'hb5c58593;
         156:    rdata = 32'h000f0517;
         157:    rdata = 32'he1850513;
         158:    rdata = 32'h6d9000ef;
         159:    rdata = 32'h4401b755;
         160:    rdata = 32'h00c4c583;
         161:    rdata = 32'h05178622;
         162:    rdata = 32'h0513000f;
         163:    rdata = 32'h10efd865;
         164:    rdata = 32'h44010ea0;
         165:    rdata = 32'h41dcb771;
         166:    rdata = 32'hc6061141;
         167:    rdata = 32'h02f04063;
         168:    rdata = 32'h00002597;
         169:    rdata = 32'hb4058593;
         170:    rdata = 32'h000f0517;
         171:    rdata = 32'hde050513;
         172:    rdata = 32'h6a1000ef;
         173:    rdata = 32'h40b24505;
         174:    rdata = 32'h80820141;
         175:    rdata = 32'h47854598;
         176:    rdata = 32'h00f70763;
         177:    rdata = 32'h00002597;
         178:    rdata = 32'hb3858593;
         179:    rdata = 32'hc583bff1;
         180:    rdata = 32'h051700c5;
         181:    rdata = 32'h0513000f;
         182:    rdata = 32'h10efd3a5;
         183:    rdata = 32'h25970b40;
         184:    rdata = 32'h85930000;
         185:    rdata = 32'hc509ae25;
         186:    rdata = 32'h00002597;
         187:    rdata = 32'had458593;
         188:    rdata = 32'h000f0517;
         189:    rdata = 32'hd9850513;
         190:    rdata = 32'h659000ef;
         191:    rdata = 32'h00002597;
         192:    rdata = 32'hb1c58593;
         193:    rdata = 32'h64d000ef;
         194:    rdata = 32'hb7754501;
         195:    rdata = 32'h114141dc;
         196:    rdata = 32'h4705c606;
         197:    rdata = 32'h02f74063;
         198:    rdata = 32'h00002597;
         199:    rdata = 32'ha6458593;
         200:    rdata = 32'h000f0517;
         201:    rdata = 32'hd6850513;
         202:    rdata = 32'h629000ef;
         203:    rdata = 32'h40b24505;
         204:    rdata = 32'h80820141;
         205:    rdata = 32'h9563459c;
         206:    rdata = 32'h519800e7;
         207:    rdata = 32'h00f70763;
         208:    rdata = 32'h00002597;
         209:    rdata = 32'ha5858593;
         210:    rdata = 32'h51d0bfe1;
         211:    rdata = 32'h00c5c583;
         212:    rdata = 32'h000f0517;
         213:    rdata = 32'hcbc50513;
         214:    rdata = 32'h00c03633;
         215:    rdata = 32'h066010ef;
         216:    rdata = 32'hb7f14501;
         217:    rdata = 32'h110141dc;
         218:    rdata = 32'h4063ce06;
         219:    rdata = 32'h259702f0;
         220:    rdata = 32'h85930000;
         221:    rdata = 32'h0517a725;
         222:    rdata = 32'h0513000f;
         223:    rdata = 32'h00efd125;
         224:    rdata = 32'h45055d30;
         225:    rdata = 32'h610540f2;
         226:    rdata = 32'h45988082;
         227:    rdata = 32'h07634785;
         228:    rdata = 32'h259700f7;
         229:    rdata = 32'h85930000;
         230:    rdata = 32'hbff1a6a5;
         231:    rdata = 32'h00c5c583;
         232:    rdata = 32'h000f0517;
         233:    rdata = 32'hc6c50513;
         234:    rdata = 32'h7f9000ef;
         235:    rdata = 32'h006cc62a;
         236:    rdata = 32'h000f0517;
         237:    rdata = 32'hcd850513;
         238:    rdata = 32'h5b5000ef;
         239:    rdata = 32'h00002597;
         240:    rdata = 32'ha5c58593;
         241:    rdata = 32'h58d000ef;
         242:    rdata = 32'hbf6d4501;
         243:    rdata = 32'h114141dc;
         244:    rdata = 32'hc422c606;
         245:    rdata = 32'h02f04163;
         246:    rdata = 32'h00002597;
         247:    rdata = 32'ha0858593;
         248:    rdata = 32'h000f0517;
         249:    rdata = 32'hca850513;
         250:    rdata = 32'h569000ef;
         251:    rdata = 32'h40b24505;
         252:    rdata = 32'h01414422;
         253:    rdata = 32'h45988082;
         254:    rdata = 32'h842e4785;
         255:    rdata = 32'h00f70763;
         256:    rdata = 32'h00002597;
         257:    rdata = 32'h9fc58593;
         258:    rdata = 32'h45dcbfe1;
         259:    rdata = 32'h04f05363;
         260:    rdata = 32'h00000597;
         261:    rdata = 32'hd8458593;
         262:    rdata = 32'h000f0517;
         263:    rdata = 32'hbe850513;
         264:    rdata = 32'h611000ef;
         265:    rdata = 32'h6731445c;
         266:    rdata = 32'h35070713;
         267:    rdata = 32'h02e787b3;
         268:    rdata = 32'h000f0517;
         269:    rdata = 32'hc3050513;
         270:    rdata = 32'h17fd4558;
         271:    rdata = 32'h10efc31c;
         272:    rdata = 32'h05171de0;
         273:    rdata = 32'h0513000f;
         274:    rdata = 32'h00efbbe5;
         275:    rdata = 32'h45015c50;
         276:    rdata = 32'h0517bf79;
         277:    rdata = 32'h0513000f;
         278:    rdata = 32'h10efc0e5;
         279:    rdata = 32'h05171ce0;
         280:    rdata = 32'h0513000f;
         281:    rdata = 32'h00efba25;
         282:    rdata = 32'hb7d55d70;
         283:    rdata = 32'h110141d8;
         284:    rdata = 32'hcc22ce06;
         285:    rdata = 32'h4789ca26;
         286:    rdata = 32'h02e7c363;
         287:    rdata = 32'h00002597;
         288:    rdata = 32'h90058593;
         289:    rdata = 32'h000f0517;
         290:    rdata = 32'hc0450513;
         291:    rdata = 32'h4c5000ef;
         292:    rdata = 32'h40f24405;
         293:    rdata = 32'h44628522;
         294:    rdata = 32'h610544d2;
         295:    rdata = 32'h459c8082;
         296:    rdata = 32'h97634705;
         297:    rdata = 32'h518000e7;
         298:    rdata = 32'h5d84e401;
         299:    rdata = 32'h00f48763;
         300:    rdata = 32'h00002597;
         301:    rdata = 32'h8e858593;
         302:    rdata = 32'hc783b7f1;
         303:    rdata = 32'h07130245;
         304:    rdata = 32'h846302d0;
         305:    rdata = 32'h666306e7;
         306:    rdata = 32'h071302f7;
         307:    rdata = 32'h826302a0;
         308:    rdata = 32'h071306e7;
         309:    rdata = 32'h886302b0;
         310:    rdata = 32'h259702e7;
         311:    rdata = 32'h85930000;
         312:    rdata = 32'h051795e5;
         313:    rdata = 32'h0513000f;
         314:    rdata = 32'h00efba65;
         315:    rdata = 32'h84264670;
         316:    rdata = 32'h0713b74d;
         317:    rdata = 32'h92e302f0;
         318:    rdata = 32'h5dd8fee7;
         319:    rdata = 32'h45dcc321;
         320:    rdata = 32'h02e7c7b3;
         321:    rdata = 32'h45dca021;
         322:    rdata = 32'h97ba5dd8;
         323:    rdata = 32'h0517006c;
         324:    rdata = 32'h0513000f;
         325:    rdata = 32'hc63eb7a5;
         326:    rdata = 32'h455000ef;
         327:    rdata = 32'h00002597;
         328:    rdata = 32'h8fc58593;
         329:    rdata = 32'h42d000ef;
         330:    rdata = 32'h45dcb7ad;
         331:    rdata = 32'h8f995dd8;
         332:    rdata = 32'h45dcbff1;
         333:    rdata = 32'h87b35dd8;
         334:    rdata = 32'hbfc902e7;
         335:    rdata = 32'h00002597;
         336:    rdata = 32'h8e058593;
         337:    rdata = 32'h1101b781;
         338:    rdata = 32'hcc22ce06;
         339:    rdata = 32'h0113ca26;
         340:    rdata = 32'h06138101;
         341:    rdata = 32'h45810400;
         342:    rdata = 32'h10ef850a;
         343:    rdata = 32'h858a2fa0;
         344:    rdata = 32'h000f0517;
         345:    rdata = 32'had050513;
         346:    rdata = 32'h739000ef;
         347:    rdata = 32'h000f0517;
         348:    rdata = 32'ha9450513;
         349:    rdata = 32'h47b000ef;
         350:    rdata = 32'h4601842a;
         351:    rdata = 32'h000f0597;
         352:    rdata = 32'hb0858593;
         353:    rdata = 32'h00ef850a;
         354:    rdata = 32'h05175cc0;
         355:    rdata = 32'h0513000f;
         356:    rdata = 32'h00efa765;
         357:    rdata = 32'h05b345d0;
         358:    rdata = 32'h25174085;
         359:    rdata = 32'h05130000;
         360:    rdata = 32'h21b98be5;
         361:    rdata = 32'h0084840a;
         362:    rdata = 32'h7c045503;
         363:    rdata = 32'h26f50409;
         364:    rdata = 32'hfe941ce3;
         365:    rdata = 32'h7f010113;
         366:    rdata = 32'h446240f2;
         367:    rdata = 32'h610544d2;
         368:    rdata = 32'h715d8082;
         369:    rdata = 32'h04000593;
         370:    rdata = 32'h000f0517;
         371:    rdata = 32'ha6850513;
         372:    rdata = 32'hc4a2c686;
         373:    rdata = 32'h6fb000ef;
         374:    rdata = 32'h04000613;
         375:    rdata = 32'h850a4581;
         376:    rdata = 32'h274010ef;
         377:    rdata = 32'h0517858a;
         378:    rdata = 32'h0513000f;
         379:    rdata = 32'h00efa4a5;
         380:    rdata = 32'h05176b30;
         381:    rdata = 32'h0513000f;
         382:    rdata = 32'h00efa0e5;
         383:    rdata = 32'h842a3f50;
         384:    rdata = 32'h000f0517;
         385:    rdata = 32'ha8450513;
         386:    rdata = 32'h6b0000ef;
         387:    rdata = 32'h000f0517;
         388:    rdata = 32'h9f450513;
         389:    rdata = 32'h3db000ef;
         390:    rdata = 32'h40850433;
         391:    rdata = 32'h00002597;
         392:    rdata = 32'h84c58593;
         393:    rdata = 32'h000f0517;
         394:    rdata = 32'ha6450513;
         395:    rdata = 32'h325000ef;
         396:    rdata = 32'h442685a2;
         397:    rdata = 32'h251740b6;
         398:    rdata = 32'h05130000;
         399:    rdata = 32'h616184e5;
         400:    rdata = 32'h712dae45;
         401:    rdata = 32'h10812c23;
         402:    rdata = 32'h10912a23;
         403:    rdata = 32'h11212823;
         404:    rdata = 32'h11312623;
         405:    rdata = 32'h11412423;
         406:    rdata = 32'h11512223;
         407:    rdata = 32'h11612023;
         408:    rdata = 32'h10112e23;
         409:    rdata = 32'h2a97842a;
         410:    rdata = 32'h8a930000;
         411:    rdata = 32'h0497832a;
         412:    rdata = 32'h8493000f;
         413:    rdata = 32'h4a2da1a4;
         414:    rdata = 32'h00001917;
         415:    rdata = 32'h36490913;
         416:    rdata = 32'h00002997;
         417:    rdata = 32'h87098993;
         418:    rdata = 32'h00002b17;
         419:    rdata = 32'h814b0b13;
         420:    rdata = 32'h852685d6;
         421:    rdata = 32'h2bd000ef;
         422:    rdata = 32'h8526004c;
         423:    rdata = 32'h279000ef;
         424:    rdata = 32'h85a20050;
         425:    rdata = 32'h24ad10a8;
         426:    rdata = 32'h63e357a6;
         427:    rdata = 32'h078afefa;
         428:    rdata = 32'h439c97ca;
         429:    rdata = 32'h878297ca;
         430:    rdata = 32'h36098522;
         431:    rdata = 32'h8522bfd1;
         432:    rdata = 32'hb7f93e01;
         433:    rdata = 32'h3e398522;
         434:    rdata = 32'h10acb7e1;
         435:    rdata = 32'h362d8522;
         436:    rdata = 32'h85ced161;
         437:    rdata = 32'ha0b18526;
         438:    rdata = 32'h852210ac;
         439:    rdata = 32'hbfcd3e6d;
         440:    rdata = 32'h852210ac;
         441:    rdata = 32'hb7ed3125;
         442:    rdata = 32'h852210ac;
         443:    rdata = 32'hb7cd39a5;
         444:    rdata = 32'h852210ac;
         445:    rdata = 32'hbfe939e1;
         446:    rdata = 32'h852210ac;
         447:    rdata = 32'hbf493b85;
         448:    rdata = 32'h35918522;
         449:    rdata = 32'h8522b771;
         450:    rdata = 32'hb7593d6d;
         451:    rdata = 32'h852685da;
         452:    rdata = 32'h241000ef;
         453:    rdata = 32'h00ef004c;
         454:    rdata = 32'h159721f0;
         455:    rdata = 32'h85930000;
         456:    rdata = 32'h00ef7a25;
         457:    rdata = 32'hb7ad22f0;
         458:    rdata = 32'h0713852e;
         459:    rdata = 32'h47830200;
         460:    rdata = 32'hc7890005;
         461:    rdata = 32'h00e79563;
         462:    rdata = 32'hbfd50505;
         463:    rdata = 32'h80824501;
         464:    rdata = 32'h00064783;
         465:    rdata = 32'h0df7f713;
         466:    rdata = 32'h0585c711;
         467:    rdata = 32'h8fa30605;
         468:    rdata = 32'hb7fdfef5;
         469:    rdata = 32'h00058023;
         470:    rdata = 32'hc7838082;
         471:    rdata = 32'hf7930005;
         472:    rdata = 32'hc3990df7;
         473:    rdata = 32'hbfd50585;
         474:    rdata = 32'hfff58513;
         475:    rdata = 32'h11018082;
         476:    rdata = 32'hc84acc22;
         477:    rdata = 32'hc256c452;
         478:    rdata = 32'hce06c05a;
         479:    rdata = 32'hc64eca26;
         480:    rdata = 32'h8432892a;
         481:    rdata = 32'h0a134b15;
         482:    rdata = 32'h4ae10086;
         483:    rdata = 32'h46634044;
         484:    rdata = 32'h854a029b;
         485:    rdata = 32'h89aa3f51;
         486:    rdata = 32'h85b3c10d;
         487:    rdata = 32'h862a0354;
         488:    rdata = 32'h0591854a;
         489:    rdata = 32'h3f6995d2;
         490:    rdata = 32'h854a85ce;
         491:    rdata = 32'h405c377d;
         492:    rdata = 32'h00150593;
         493:    rdata = 32'hc05c0785;
         494:    rdata = 32'h40f2bfd1;
         495:    rdata = 32'h44d24462;
         496:    rdata = 32'h49b24942;
         497:    rdata = 32'h4a924a22;
         498:    rdata = 32'h61054b02;
         499:    rdata = 32'h11418082;
         500:    rdata = 32'h8493c226;
         501:    rdata = 32'hc42200c5;
         502:    rdata = 32'h842e8526;
         503:    rdata = 32'h00001597;
         504:    rdata = 32'h72c58593;
         505:    rdata = 32'h00efc606;
         506:    rdata = 32'he9197020;
         507:    rdata = 32'h00042023;
         508:    rdata = 32'h40b2405c;
         509:    rdata = 32'h17fd4492;
         510:    rdata = 32'h4422c05c;
         511:    rdata = 32'h80820141;
         512:    rdata = 32'h00001597;
         513:    rdata = 32'h71058593;
         514:    rdata = 32'h00ef8526;
         515:    rdata = 32'h47856de0;
         516:    rdata = 32'h1597c14d;
         517:    rdata = 32'h85930000;
         518:    rdata = 32'h85267065;
         519:    rdata = 32'h6cc000ef;
         520:    rdata = 32'hc9414789;
         521:    rdata = 32'h00001597;
         522:    rdata = 32'h6fc58593;
         523:    rdata = 32'h00ef8526;
         524:    rdata = 32'h478d6ba0;
         525:    rdata = 32'h1597cd3d;
         526:    rdata = 32'h85930000;
         527:    rdata = 32'h85266fe5;
         528:    rdata = 32'h6a8000ef;
         529:    rdata = 32'hc5354791;
         530:    rdata = 32'h00001597;
         531:    rdata = 32'h70058593;
         532:    rdata = 32'h00ef8526;
         533:    rdata = 32'h47956960;
         534:    rdata = 32'h1597cd29;
         535:    rdata = 32'h85930000;
         536:    rdata = 32'h85266fa5;
         537:    rdata = 32'h684000ef;
         538:    rdata = 32'hc5214799;
         539:    rdata = 32'h00001597;
         540:    rdata = 32'h6f458593;
         541:    rdata = 32'h00ef8526;
         542:    rdata = 32'h479d6720;
         543:    rdata = 32'h1597c91d;
         544:    rdata = 32'h85930000;
         545:    rdata = 32'h85266f25;
         546:    rdata = 32'h660000ef;
         547:    rdata = 32'hc11547a1;
         548:    rdata = 32'h00001597;
         549:    rdata = 32'h6ec58593;
         550:    rdata = 32'h25b98526;
         551:    rdata = 32'hc91147a5;
         552:    rdata = 32'h00001597;
         553:    rdata = 32'h6e858593;
         554:    rdata = 32'h2d3d8526;
         555:    rdata = 32'hc11147a9;
         556:    rdata = 32'hc01c47ad;
         557:    rdata = 32'h1101bf35;
         558:    rdata = 32'hc84acc22;
         559:    rdata = 32'hc452c64e;
         560:    rdata = 32'hca26ce06;
         561:    rdata = 32'h8413892e;
         562:    rdata = 32'h498100c5;
         563:    rdata = 32'h27834a05;
         564:    rdata = 32'hd7630049;
         565:    rdata = 32'h049302f9;
         566:    rdata = 32'h85260184;
         567:    rdata = 32'h00ef0985;
         568:    rdata = 32'hc9097420;
         569:    rdata = 32'hff442e23;
         570:    rdata = 32'h00ef8526;
         571:    rdata = 32'hc00876c0;
         572:    rdata = 32'hbff18426;
         573:    rdata = 32'hfe042e23;
         574:    rdata = 32'h852285a6;
         575:    rdata = 32'hbfcd2b7d;
         576:    rdata = 32'h446240f2;
         577:    rdata = 32'h494244d2;
         578:    rdata = 32'h4a2249b2;
         579:    rdata = 32'h80826105;
         580:    rdata = 32'hc6061141;
         581:    rdata = 32'hc226c422;
         582:    rdata = 32'h842ac04a;
         583:    rdata = 32'h893284ae;
         584:    rdata = 32'h00052223;
         585:    rdata = 32'h09000613;
         586:    rdata = 32'h05214581;
         587:    rdata = 32'h729000ef;
         588:    rdata = 32'h85ca8622;
         589:    rdata = 32'h3d258526;
         590:    rdata = 32'heb91405c;
         591:    rdata = 32'hc01c47b1;
         592:    rdata = 32'h852240b2;
         593:    rdata = 32'h44924422;
         594:    rdata = 32'h01414902;
         595:    rdata = 32'h85a28082;
         596:    rdata = 32'h3db58526;
         597:    rdata = 32'h852685a2;
         598:    rdata = 32'hb7dd3fb9;
         599:    rdata = 32'h85aa7119;
         600:    rdata = 32'hde860068;
         601:    rdata = 32'h15972b99;
         602:    rdata = 32'h85930000;
         603:    rdata = 32'h00684b25;
         604:    rdata = 32'h006c2bb1;
         605:    rdata = 32'h000ef517;
         606:    rdata = 32'h71450513;
         607:    rdata = 32'h7d4000ef;
         608:    rdata = 32'h610950f6;
         609:    rdata = 32'h11018082;
         610:    rdata = 32'h004885aa;
         611:    rdata = 32'h23ddce06;
         612:    rdata = 32'h37e90048;
         613:    rdata = 32'h610540f2;
         614:    rdata = 32'h11018082;
         615:    rdata = 32'h004885aa;
         616:    rdata = 32'h2d25ce06;
         617:    rdata = 32'h3f5d0048;
         618:    rdata = 32'h610540f2;
         619:    rdata = 32'h71198082;
         620:    rdata = 32'h842edca2;
         621:    rdata = 32'h006885aa;
         622:    rdata = 32'h2301de86;
         623:    rdata = 32'h00001597;
         624:    rdata = 32'h60058593;
         625:    rdata = 32'h23190068;
         626:    rdata = 32'h006885a2;
         627:    rdata = 32'h15972301;
         628:    rdata = 32'h85930000;
         629:    rdata = 32'h006844a5;
         630:    rdata = 32'h006c29d5;
         631:    rdata = 32'h000ef517;
         632:    rdata = 32'h6ac50513;
         633:    rdata = 32'h76c000ef;
         634:    rdata = 32'h546650f6;
         635:    rdata = 32'h80826109;
         636:    rdata = 32'hcc221101;
         637:    rdata = 32'h0048842a;
         638:    rdata = 32'h2badce06;
         639:    rdata = 32'h8522004c;
         640:    rdata = 32'h40f2377d;
         641:    rdata = 32'h61054462;
         642:    rdata = 32'h11018082;
         643:    rdata = 32'h842acc22;
         644:    rdata = 32'hce060048;
         645:    rdata = 32'h004c23d9;
         646:    rdata = 32'h3f518522;
         647:    rdata = 32'h446240f2;
         648:    rdata = 32'h80826105;
         649:    rdata = 32'hdaa67119;
         650:    rdata = 32'h85aa84ae;
         651:    rdata = 32'hde860068;
         652:    rdata = 32'h8432dca2;
         653:    rdata = 32'h15972159;
         654:    rdata = 32'h85930000;
         655:    rdata = 32'h006858a5;
         656:    rdata = 32'h85a62171;
         657:    rdata = 32'h21590068;
         658:    rdata = 32'h00001597;
         659:    rdata = 32'h57c58593;
         660:    rdata = 32'h29ad0068;
         661:    rdata = 32'h006885a2;
         662:    rdata = 32'h15972995;
         663:    rdata = 32'h85930000;
         664:    rdata = 32'h00683be5;
         665:    rdata = 32'h006c21a5;
         666:    rdata = 32'h000ef517;
         667:    rdata = 32'h62050513;
         668:    rdata = 32'h6e0000ef;
         669:    rdata = 32'h546650f6;
         670:    rdata = 32'h610954d6;
         671:    rdata = 32'h71798082;
         672:    rdata = 32'h842ad422;
         673:    rdata = 32'hd6060028;
         674:    rdata = 32'h84b2d226;
         675:    rdata = 32'h85a623b9;
         676:    rdata = 32'h21cd0848;
         677:    rdata = 32'h002c0850;
         678:    rdata = 32'h37698522;
         679:    rdata = 32'h542250b2;
         680:    rdata = 32'h61455492;
         681:    rdata = 32'h71798082;
         682:    rdata = 32'h842ad422;
         683:    rdata = 32'hd6060028;
         684:    rdata = 32'h84b2d226;
         685:    rdata = 32'h85a6231d;
         686:    rdata = 32'h23050848;
         687:    rdata = 32'h002c0850;
         688:    rdata = 32'h378d8522;
         689:    rdata = 32'h542250b2;
         690:    rdata = 32'h61455492;
         691:    rdata = 32'h11018082;
         692:    rdata = 32'hce06cc22;
         693:    rdata = 32'hc84aca26;
         694:    rdata = 32'hc452c64e;
         695:    rdata = 32'h4581842a;
         696:    rdata = 32'h4585c211;
         697:    rdata = 32'h000ef517;
         698:    rdata = 32'h56c50513;
         699:    rdata = 32'h2eb000ef;
         700:    rdata = 32'h000ef517;
         701:    rdata = 32'h56050513;
         702:    rdata = 32'h201000ef;
         703:    rdata = 32'h000ef497;
         704:    rdata = 32'h55448493;
         705:    rdata = 32'h00ef8526;
         706:    rdata = 32'hdd6d1ff0;
         707:    rdata = 32'hf91744fd;
         708:    rdata = 32'h0913000e;
         709:    rdata = 32'hfa175429;
         710:    rdata = 32'h0a13000e;
         711:    rdata = 32'h59fd51aa;
         712:    rdata = 32'h00ef854a;
         713:    rdata = 32'h854a1d70;
         714:    rdata = 32'h1dd000ef;
         715:    rdata = 32'h9593dd6d;
         716:    rdata = 32'h95a20064;
         717:    rdata = 32'h14fd8552;
         718:    rdata = 32'h171000ef;
         719:    rdata = 32'hff3492e3;
         720:    rdata = 32'h852240f2;
         721:    rdata = 32'h44d24462;
         722:    rdata = 32'h49b24942;
         723:    rdata = 32'h61054a22;
         724:    rdata = 32'h11018082;
         725:    rdata = 32'h842acc22;
         726:    rdata = 32'h000ef517;
         727:    rdata = 32'h4f850513;
         728:    rdata = 32'hc62ece06;
         729:    rdata = 32'h00efc432;
         730:    rdata = 32'hf5172970;
         731:    rdata = 32'h0513000e;
         732:    rdata = 32'h00ef4e65;
         733:    rdata = 32'h46221870;
         734:    rdata = 32'h852245b2;
         735:    rdata = 32'h40f23f89;
         736:    rdata = 32'h44628522;
         737:    rdata = 32'h80826105;
         738:    rdata = 32'h878a715d;
         739:    rdata = 32'hc686c4a2;
         740:    rdata = 32'hc2a6842e;
         741:    rdata = 32'h902385be;
         742:    rdata = 32'h009800c7;
         743:    rdata = 32'h9ce30789;
         744:    rdata = 32'hf517fee7;
         745:    rdata = 32'h0513000e;
         746:    rdata = 32'h00ef48e5;
         747:    rdata = 32'h45810f70;
         748:    rdata = 32'h4585c011;
         749:    rdata = 32'h000ef517;
         750:    rdata = 32'h49c50513;
         751:    rdata = 32'h21b000ef;
         752:    rdata = 32'h000ef517;
         753:    rdata = 32'h49050513;
         754:    rdata = 32'h131000ef;
         755:    rdata = 32'h000ef417;
         756:    rdata = 32'h48440413;
         757:    rdata = 32'h00ef8522;
         758:    rdata = 32'hdd6d12f0;
         759:    rdata = 32'h02000413;
         760:    rdata = 32'h000ef497;
         761:    rdata = 32'h47048493;
         762:    rdata = 32'h00ef8526;
         763:    rdata = 32'h852610f0;
         764:    rdata = 32'h115000ef;
         765:    rdata = 32'h147ddd6d;
         766:    rdata = 32'h40b6f865;
         767:    rdata = 32'h44964426;
         768:    rdata = 32'h80826161;
         769:    rdata = 32'hca261101;
         770:    rdata = 32'hcc22ce06;
         771:    rdata = 32'hc64ec84a;
         772:    rdata = 32'he5ad84b2;
         773:    rdata = 32'h000ef517;
         774:    rdata = 32'h43c50513;
         775:    rdata = 32'h1bb000ef;
         776:    rdata = 32'h000ef517;
         777:    rdata = 32'h43050513;
         778:    rdata = 32'h0d1000ef;
         779:    rdata = 32'h000ef417;
         780:    rdata = 32'h42440413;
         781:    rdata = 32'h00ef8522;
         782:    rdata = 32'hdd6d0cf0;
         783:    rdata = 32'h7c048413;
         784:    rdata = 32'h000ef997;
         785:    rdata = 32'h3f098993;
         786:    rdata = 32'h000ef917;
         787:    rdata = 32'h40890913;
         788:    rdata = 32'h85a2854e;
         789:    rdata = 32'h04d000ef;
         790:    rdata = 32'h00ef854a;
         791:    rdata = 32'h854a09f0;
         792:    rdata = 32'h0a5000ef;
         793:    rdata = 32'h0793dd6d;
         794:    rdata = 32'h9b63fc04;
         795:    rdata = 32'h40f20084;
         796:    rdata = 32'h44d24462;
         797:    rdata = 32'h49b24942;
         798:    rdata = 32'h80826105;
         799:    rdata = 32'hbf594585;
         800:    rdata = 32'hb7f9843e;
         801:    rdata = 32'hf5171141;
         802:    rdata = 32'h0513000e;
         803:    rdata = 32'hc6063ca5;
         804:    rdata = 32'h161000ef;
         805:    rdata = 32'hf51740b2;
         806:    rdata = 32'h0513000e;
         807:    rdata = 32'h01413ba5;
         808:    rdata = 32'h0590006f;
         809:    rdata = 32'hc4221141;
         810:    rdata = 32'h842ac606;
         811:    rdata = 32'h85223fa1;
         812:    rdata = 32'h40b24422;
         813:    rdata = 32'hb7f90141;
         814:    rdata = 32'h71797379;
         815:    rdata = 32'h80030313;
         816:    rdata = 32'hd226d422;
         817:    rdata = 32'hce4ed04a;
         818:    rdata = 32'hc85acc52;
         819:    rdata = 32'hca56d606;
         820:    rdata = 32'h911a6a0d;
         821:    rdata = 32'h74fd0818;
         822:    rdata = 32'h800a0793;
         823:    rdata = 32'h849397ba;
         824:    rdata = 32'h94be8004;
         825:    rdata = 32'h842a6909;
         826:    rdata = 32'h80090613;
         827:    rdata = 32'h85264581;
         828:    rdata = 32'h365000ef;
         829:    rdata = 32'h800a0793;
         830:    rdata = 32'h97ba0818;
         831:    rdata = 32'h412787b3;
         832:    rdata = 32'hc63e4981;
         833:    rdata = 32'h02000b13;
         834:    rdata = 32'hca334901;
         835:    rdata = 32'h86520809;
         836:    rdata = 32'h85224581;
         837:    rdata = 32'h45853d95;
         838:    rdata = 32'h4ab38522;
         839:    rdata = 32'h86560809;
         840:    rdata = 32'h852235a5;
         841:    rdata = 32'h45323785;
         842:    rdata = 32'h85a24601;
         843:    rdata = 32'h4732351d;
         844:    rdata = 32'h86ba87a6;
         845:    rdata = 32'h0c078593;
         846:    rdata = 32'h0006d603;
         847:    rdata = 32'h0047d503;
         848:    rdata = 32'h00c57863;
         849:    rdata = 32'h01479023;
         850:    rdata = 32'h01579123;
         851:    rdata = 32'h00c79223;
         852:    rdata = 32'h06890799;
         853:    rdata = 32'hfeb792e3;
         854:    rdata = 32'h8693668d;
         855:    rdata = 32'h08108006;
         856:    rdata = 32'h071396b2;
         857:    rdata = 32'h96e30407;
         858:    rdata = 32'h0905fcf6;
         859:    rdata = 32'hfb6911e3;
         860:    rdata = 32'h9be30985;
         861:    rdata = 32'h660df929;
         862:    rdata = 32'h80060713;
         863:    rdata = 32'h05130814;
         864:    rdata = 32'h08048006;
         865:    rdata = 32'h80060613;
         866:    rdata = 32'h77fd9736;
         867:    rdata = 32'h962676f9;
         868:    rdata = 32'h859397ba;
         869:    rdata = 32'h95268006;
         870:    rdata = 32'h95aa96b2;
         871:    rdata = 32'h80278793;
         872:    rdata = 32'hc6364701;
         873:    rdata = 32'h04000513;
         874:    rdata = 32'h8e3346b2;
         875:    rdata = 32'h863e00e5;
         876:    rdata = 32'h00e68333;
         877:    rdata = 32'h58834681;
         878:    rdata = 32'h0833ffe6;
         879:    rdata = 32'h061900de;
         880:    rdata = 32'h01181023;
         881:    rdata = 32'hffa65883;
         882:    rdata = 32'h00d30833;
         883:    rdata = 32'h10230689;
         884:    rdata = 32'h92e30118;
         885:    rdata = 32'h0713fea6;
         886:    rdata = 32'h06930407;
         887:    rdata = 32'h87938007;
         888:    rdata = 32'hf2f90c07;
         889:    rdata = 32'h0818690d;
         890:    rdata = 32'h079374f9;
         891:    rdata = 32'h97ba8009;
         892:    rdata = 32'h80048613;
         893:    rdata = 32'h8522963e;
         894:    rdata = 32'h356d4581;
         895:    rdata = 32'h07930818;
         896:    rdata = 32'h97ba8009;
         897:    rdata = 32'h00978633;
         898:    rdata = 32'h45858522;
         899:    rdata = 32'h630d3d61;
         900:    rdata = 32'h80030313;
         901:    rdata = 32'h50b2911a;
         902:    rdata = 32'h54925422;
         903:    rdata = 32'h49f25902;
         904:    rdata = 32'h4ad24a62;
         905:    rdata = 32'h61454b42;
         906:    rdata = 32'h11418082;
         907:    rdata = 32'hc606c422;
         908:    rdata = 32'h3b99842a;
         909:    rdata = 32'h44228522;
         910:    rdata = 32'h014140b2;
         911:    rdata = 32'h0713b5a1;
         912:    rdata = 32'h47830300;
         913:    rdata = 32'h94630005;
         914:    rdata = 32'h050500e7;
         915:    rdata = 32'he391bfdd;
         916:    rdata = 32'h8082157d;
         917:    rdata = 32'h00054703;
         918:    rdata = 32'h02d00793;
         919:    rdata = 32'h00f71363;
         920:    rdata = 32'h47250505;
         921:    rdata = 32'h00054783;
         922:    rdata = 32'hfd078793;
         923:    rdata = 32'h0ff7f793;
         924:    rdata = 32'h00f76863;
         925:    rdata = 32'h00154783;
         926:    rdata = 32'hf7ed0505;
         927:    rdata = 32'h80824505;
         928:    rdata = 32'h80824501;
         929:    rdata = 32'h46a50509;
         930:    rdata = 32'h47834615;
         931:    rdata = 32'h87130005;
         932:    rdata = 32'h7713fd07;
         933:    rdata = 32'hfa630ff7;
         934:    rdata = 32'hf79300e6;
         935:    rdata = 32'h8793fdf7;
         936:    rdata = 32'hf793fbf7;
         937:    rdata = 32'h68630ff7;
         938:    rdata = 32'h478300f6;
         939:    rdata = 32'h05050015;
         940:    rdata = 32'h4505ffe9;
         941:    rdata = 32'h45018082;
         942:    rdata = 32'h87aa8082;
         943:    rdata = 32'h0005c703;
         944:    rdata = 32'h07850585;
         945:    rdata = 32'hfee78fa3;
         946:    rdata = 32'h8082fb75;
         947:    rdata = 32'hc68387aa;
         948:    rdata = 32'h873e0007;
         949:    rdata = 32'hfee50785;
         950:    rdata = 32'h0005c783;
         951:    rdata = 32'h07050585;
         952:    rdata = 32'hfef70fa3;
         953:    rdata = 32'h8082fbf5;
         954:    rdata = 32'h00054783;
         955:    rdata = 32'h0005c703;
         956:    rdata = 32'h00e78763;
         957:    rdata = 32'he963557d;
         958:    rdata = 32'h450500e7;
         959:    rdata = 32'hc7818082;
         960:    rdata = 32'h05850505;
         961:    rdata = 32'h4501b7d5;
         962:    rdata = 32'h87aa8082;
         963:    rdata = 32'h87334501;
         964:    rdata = 32'h470300a7;
         965:    rdata = 32'hc3190007;
         966:    rdata = 32'hbfd50505;
         967:    rdata = 32'h47898082;
         968:    rdata = 32'h02f60c63;
         969:    rdata = 32'h0d634791;
         970:    rdata = 32'h470502f6;
         971:    rdata = 32'h14634781;
         972:    rdata = 32'h079300e6;
         973:    rdata = 32'h46290640;
         974:    rdata = 32'hd733cb8d;
         975:    rdata = 32'h050502f5;
         976:    rdata = 32'h0ff77693;
         977:    rdata = 32'h02f686b3;
         978:    rdata = 32'h03070713;
         979:    rdata = 32'hfee50fa3;
         980:    rdata = 32'h02c7d7b3;
         981:    rdata = 32'hb7cd8d95;
         982:    rdata = 32'h87936789;
         983:    rdata = 32'hbfe17107;
         984:    rdata = 32'h3b9ad7b7;
         985:    rdata = 32'ha0078793;
         986:    rdata = 32'h0023b7f9;
         987:    rdata = 32'h80820005;
         988:    rdata = 32'hb7754605;
         989:    rdata = 32'hcc221101;
         990:    rdata = 32'h842a4611;
         991:    rdata = 32'hce060048;
         992:    rdata = 32'h00483f79;
         993:    rdata = 32'h85aa3d6d;
         994:    rdata = 32'h3f058522;
         995:    rdata = 32'h446240f2;
         996:    rdata = 32'h80826105;
         997:    rdata = 32'h03000793;
         998:    rdata = 32'h76130606;
         999:    rdata = 32'h00230ff6;
        1000:    rdata = 32'h079300f5;
        1001:    rdata = 32'h00a30780;
        1002:    rdata = 32'h482500f5;
        1003:    rdata = 32'hc38587b2;
        1004:    rdata = 32'h00f5f713;
        1005:    rdata = 32'h05770693;
        1006:    rdata = 32'h00e86463;
        1007:    rdata = 32'h03070693;
        1008:    rdata = 32'h00f50733;
        1009:    rdata = 32'h00d700a3;
        1010:    rdata = 32'h17fd8191;
        1011:    rdata = 32'h9532b7cd;
        1012:    rdata = 32'h00050123;
        1013:    rdata = 32'h46058082;
        1014:    rdata = 32'h4611bf75;
        1015:    rdata = 32'h1101bf65;
        1016:    rdata = 32'hce06cc22;
        1017:    rdata = 32'hd563842a;
        1018:    rdata = 32'h07130205;
        1019:    rdata = 32'h002302d0;
        1020:    rdata = 32'h05b300e5;
        1021:    rdata = 32'h461140b0;
        1022:    rdata = 32'h37150048;
        1023:    rdata = 32'h35810048;
        1024:    rdata = 32'h051385aa;
        1025:    rdata = 32'h3d550014;
        1026:    rdata = 32'h446240f2;
        1027:    rdata = 32'h80826105;
        1028:    rdata = 32'h00484611;
        1029:    rdata = 32'h00483729;
        1030:    rdata = 32'h85aa351d;
        1031:    rdata = 32'hb7e58522;
        1032:    rdata = 32'hc4221141;
        1033:    rdata = 32'h842ac606;
        1034:    rdata = 32'he1153535;
        1035:    rdata = 32'h00044703;
        1036:    rdata = 32'h03000793;
        1037:    rdata = 32'h00f71d63;
        1038:    rdata = 32'h00144703;
        1039:    rdata = 32'h07800793;
        1040:    rdata = 32'h00f71763;
        1041:    rdata = 32'h44228522;
        1042:    rdata = 32'h014140b2;
        1043:    rdata = 32'h40b2bd25;
        1044:    rdata = 32'h01414422;
        1045:    rdata = 32'h11418082;
        1046:    rdata = 32'hc606c422;
        1047:    rdata = 32'h3bdd842a;
        1048:    rdata = 32'h00044783;
        1049:    rdata = 32'h0693c91d;
        1050:    rdata = 32'h470102d0;
        1051:    rdata = 32'h00d79463;
        1052:    rdata = 32'h0405872a;
        1053:    rdata = 32'h46294501;
        1054:    rdata = 32'h00044683;
        1055:    rdata = 32'h07b3ca81;
        1056:    rdata = 32'h851302c5;
        1057:    rdata = 32'h0405fd06;
        1058:    rdata = 32'hb7fd953e;
        1059:    rdata = 32'h0533c319;
        1060:    rdata = 32'h40b240a0;
        1061:    rdata = 32'h01414422;
        1062:    rdata = 32'h07138082;
        1063:    rdata = 32'h96630300;
        1064:    rdata = 32'h470304e7;
        1065:    rdata = 32'h07930014;
        1066:    rdata = 32'h10630780;
        1067:    rdata = 32'h852204f7;
        1068:    rdata = 32'hcd053bd1;
        1069:    rdata = 32'h45010409;
        1070:    rdata = 32'h06000713;
        1071:    rdata = 32'h04000693;
        1072:    rdata = 32'h00044783;
        1073:    rdata = 32'h7a63d7f9;
        1074:    rdata = 32'h879300f7;
        1075:    rdata = 32'hf793fa97;
        1076:    rdata = 32'h05120ff7;
        1077:    rdata = 32'h04058d5d;
        1078:    rdata = 32'hf563b7e5;
        1079:    rdata = 32'h879300f6;
        1080:    rdata = 32'hb7f5fc97;
        1081:    rdata = 32'hfd078793;
        1082:    rdata = 32'hc537b7dd;
        1083:    rdata = 32'h0513dead;
        1084:    rdata = 32'hb745eef5;
        1085:    rdata = 32'hfdf57793;
        1086:    rdata = 32'hfbf78793;
        1087:    rdata = 32'h0ff7f793;
        1088:    rdata = 32'h77634765;
        1089:    rdata = 32'h051300f7;
        1090:    rdata = 32'h3513fd05;
        1091:    rdata = 32'h808200a5;
        1092:    rdata = 32'h80824505;
        1093:    rdata = 32'hc4221141;
        1094:    rdata = 32'h06400613;
        1095:    rdata = 32'hf517842a;
        1096:    rdata = 32'h0513000e;
        1097:    rdata = 32'hc606f525;
        1098:    rdata = 32'h40b22b89;
        1099:    rdata = 32'h44228522;
        1100:    rdata = 32'h80820141;
        1101:    rdata = 32'hc4221141;
        1102:    rdata = 32'hf517842a;
        1103:    rdata = 32'h0513000e;
        1104:    rdata = 32'hc606f365;
        1105:    rdata = 32'h40b22365;
        1106:    rdata = 32'h44228522;
        1107:    rdata = 32'h80820141;
        1108:    rdata = 32'hc4221141;
        1109:    rdata = 32'hf517842a;
        1110:    rdata = 32'h0513000e;
        1111:    rdata = 32'hc606f1a5;
        1112:    rdata = 32'h40b22371;
        1113:    rdata = 32'h44228522;
        1114:    rdata = 32'h80820141;
        1115:    rdata = 32'h1101418c;
        1116:    rdata = 32'h842acc22;
        1117:    rdata = 32'hce060048;
        1118:    rdata = 32'h004c359d;
        1119:    rdata = 32'h000ef517;
        1120:    rdata = 32'hef450513;
        1121:    rdata = 32'h40f223a5;
        1122:    rdata = 32'h44628522;
        1123:    rdata = 32'h80826105;
        1124:    rdata = 32'hc5227175;
        1125:    rdata = 32'hc14ac326;
        1126:    rdata = 32'hdcd2dece;
        1127:    rdata = 32'h84aac706;
        1128:    rdata = 32'hf417892e;
        1129:    rdata = 32'h0413000e;
        1130:    rdata = 32'h1a17ece4;
        1131:    rdata = 32'h0a130000;
        1132:    rdata = 32'h1997e12a;
        1133:    rdata = 32'h89930000;
        1134:    rdata = 32'h85cae169;
        1135:    rdata = 32'h233d8522;
        1136:    rdata = 32'h852285d2;
        1137:    rdata = 32'h006c2325;
        1138:    rdata = 32'h37a98526;
        1139:    rdata = 32'h3d890068;
        1140:    rdata = 32'h85cee509;
        1141:    rdata = 32'h2b198522;
        1142:    rdata = 32'h0068b7cd;
        1143:    rdata = 32'h40ba3dad;
        1144:    rdata = 32'h449a442a;
        1145:    rdata = 32'h59f6490a;
        1146:    rdata = 32'h61495a66;
        1147:    rdata = 32'h25738082;
        1148:    rdata = 32'h25f3b000;
        1149:    rdata = 32'h8082b800;
        1150:    rdata = 32'h00010001;
        1151:    rdata = 32'h00010001;
        1152:    rdata = 32'h00010001;
        1153:    rdata = 32'hf9ed15fd;
        1154:    rdata = 32'hc10c8082;
        1155:    rdata = 32'h62f38082;
        1156:    rdata = 32'h80823004;
        1157:    rdata = 32'h300472f3;
        1158:    rdata = 32'hc14c8082;
        1159:    rdata = 32'ha2f362c1;
        1160:    rdata = 32'h80823042;
        1161:    rdata = 32'h00052223;
        1162:    rdata = 32'hb2f362c1;
        1163:    rdata = 32'h80823042;
        1164:    rdata = 32'h02b7c50c;
        1165:    rdata = 32'ha2f30002;
        1166:    rdata = 32'h80823042;
        1167:    rdata = 32'h00052423;
        1168:    rdata = 32'h000202b7;
        1169:    rdata = 32'h3042b2f3;
        1170:    rdata = 32'h71398082;
        1171:    rdata = 32'hde06cc3e;
        1172:    rdata = 32'hda1adc16;
        1173:    rdata = 32'hd62ad81e;
        1174:    rdata = 32'hd232d42e;
        1175:    rdata = 32'hce3ad036;
        1176:    rdata = 32'hc846ca42;
        1177:    rdata = 32'hc476c672;
        1178:    rdata = 32'hc07ec27a;
        1179:    rdata = 32'h000ef797;
        1180:    rdata = 32'hd947a783;
        1181:    rdata = 32'h9782c78d;
        1182:    rdata = 32'h52e250f2;
        1183:    rdata = 32'h53c25352;
        1184:    rdata = 32'h55a25532;
        1185:    rdata = 32'h56825612;
        1186:    rdata = 32'h47e24772;
        1187:    rdata = 32'h48c24852;
        1188:    rdata = 32'h4ea24e32;
        1189:    rdata = 32'h4f824f12;
        1190:    rdata = 32'h00736121;
        1191:    rdata = 32'ha0013020;
        1192:    rdata = 32'hcc3e7139;
        1193:    rdata = 32'hdc16de06;
        1194:    rdata = 32'hd81eda1a;
        1195:    rdata = 32'hd42ed62a;
        1196:    rdata = 32'hd036d232;
        1197:    rdata = 32'hca42ce3a;
        1198:    rdata = 32'hc672c846;
        1199:    rdata = 32'hc27ac476;
        1200:    rdata = 32'hf797c07e;
        1201:    rdata = 32'ha783000e;
        1202:    rdata = 32'h9782d427;
        1203:    rdata = 32'h52e250f2;
        1204:    rdata = 32'h53c25352;
        1205:    rdata = 32'h55a25532;
        1206:    rdata = 32'h56825612;
        1207:    rdata = 32'h47e24772;
        1208:    rdata = 32'h48c24852;
        1209:    rdata = 32'h4ea24e32;
        1210:    rdata = 32'h4f824f12;
        1211:    rdata = 32'h00736121;
        1212:    rdata = 32'h71393020;
        1213:    rdata = 32'hde06cc3e;
        1214:    rdata = 32'hda1adc16;
        1215:    rdata = 32'hd62ad81e;
        1216:    rdata = 32'hd232d42e;
        1217:    rdata = 32'hce3ad036;
        1218:    rdata = 32'hc846ca42;
        1219:    rdata = 32'hc476c672;
        1220:    rdata = 32'hc07ec27a;
        1221:    rdata = 32'h000ef797;
        1222:    rdata = 32'hcf47a783;
        1223:    rdata = 32'h50f29782;
        1224:    rdata = 32'h535252e2;
        1225:    rdata = 32'h553253c2;
        1226:    rdata = 32'h561255a2;
        1227:    rdata = 32'h47725682;
        1228:    rdata = 32'h485247e2;
        1229:    rdata = 32'h4e3248c2;
        1230:    rdata = 32'h4f124ea2;
        1231:    rdata = 32'h61214f82;
        1232:    rdata = 32'h30200073;
        1233:    rdata = 32'h00458793;
        1234:    rdata = 32'h8793c15c;
        1235:    rdata = 32'hc51c0085;
        1236:    rdata = 32'h00c58793;
        1237:    rdata = 32'h8793c55c;
        1238:    rdata = 32'hc91c0105;
        1239:    rdata = 32'h01458793;
        1240:    rdata = 32'h8793c95c;
        1241:    rdata = 32'hc10c0185;
        1242:    rdata = 32'h8793cd1c;
        1243:    rdata = 32'h859301c5;
        1244:    rdata = 32'hcd5c0205;
        1245:    rdata = 32'h8082d10c;
        1246:    rdata = 32'h8a05511c;
        1247:    rdata = 32'h00b61633;
        1248:    rdata = 32'h97b3439c;
        1249:    rdata = 32'h8e5d48b7;
        1250:    rdata = 32'hc390511c;
        1251:    rdata = 32'h511c8082;
        1252:    rdata = 32'h47854388;
        1253:    rdata = 32'h00b797b3;
        1254:    rdata = 32'h35338d7d;
        1255:    rdata = 32'h808200a0;
        1256:    rdata = 32'h4388455c;
        1257:    rdata = 32'h97b34785;
        1258:    rdata = 32'h8d7d00b7;
        1259:    rdata = 32'h00a03533;
        1260:    rdata = 32'h451c8082;
        1261:    rdata = 32'h8e3d439c;
        1262:    rdata = 32'h8e3d8e6d;
        1263:    rdata = 32'hc390451c;
        1264:    rdata = 32'h47858082;
        1265:    rdata = 32'h00b61633;
        1266:    rdata = 32'h00b795b3;
        1267:    rdata = 32'h1141b7dd;
        1268:    rdata = 32'hc226c422;
        1269:    rdata = 32'h842ac606;
        1270:    rdata = 32'h37d984ae;
        1271:    rdata = 32'h00154613;
        1272:    rdata = 32'h44228522;
        1273:    rdata = 32'h85a640b2;
        1274:    rdata = 32'h76134492;
        1275:    rdata = 32'h01410ff6;
        1276:    rdata = 32'h455cbfc9;
        1277:    rdata = 32'h55134388;
        1278:    rdata = 32'h80824915;
        1279:    rdata = 32'h4388455c;
        1280:    rdata = 32'h49055513;
        1281:    rdata = 32'h11418082;
        1282:    rdata = 32'h4601c226;
        1283:    rdata = 32'h45bd84ae;
        1284:    rdata = 32'hc606c422;
        1285:    rdata = 32'h378d842a;
        1286:    rdata = 32'h44228522;
        1287:    rdata = 32'h862640b2;
        1288:    rdata = 32'h45bd4492;
        1289:    rdata = 32'hbf710141;
        1290:    rdata = 32'h00858713;
        1291:    rdata = 32'h8793c518;
        1292:    rdata = 32'h87130505;
        1293:    rdata = 32'hc55800c5;
        1294:    rdata = 32'h8713c95c;
        1295:    rdata = 32'h07b70105;
        1296:    rdata = 32'hc9180101;
        1297:    rdata = 32'h00458613;
        1298:    rdata = 32'h10078713;
        1299:    rdata = 32'h20078793;
        1300:    rdata = 32'hc150c10c;
        1301:    rdata = 32'hcd5ccd18;
        1302:    rdata = 32'h02050513;
        1303:    rdata = 32'h4118a8a5;
        1304:    rdata = 32'h97938985;
        1305:    rdata = 32'h430c0025;
        1306:    rdata = 32'h8ddd99ed;
        1307:    rdata = 32'h8082c30c;
        1308:    rdata = 32'h89854118;
        1309:    rdata = 32'h00359793;
        1310:    rdata = 32'h99dd430c;
        1311:    rdata = 32'hc30c8ddd;
        1312:    rdata = 32'h41188082;
        1313:    rdata = 32'h97938985;
        1314:    rdata = 32'h430c0045;
        1315:    rdata = 32'h8ddd99bd;
        1316:    rdata = 32'h8082c30c;
        1317:    rdata = 32'hc38c451c;
        1318:    rdata = 32'h455c8082;
        1319:    rdata = 32'h80824388;
        1320:    rdata = 32'h06134908;
        1321:    rdata = 32'hac490400;
        1322:    rdata = 32'h852e87aa;
        1323:    rdata = 32'h06134bcc;
        1324:    rdata = 32'ha4590400;
        1325:    rdata = 32'h41984d1c;
        1326:    rdata = 32'h4d1cc398;
        1327:    rdata = 32'hc3d841d8;
        1328:    rdata = 32'h4d1c4598;
        1329:    rdata = 32'h45d8c798;
        1330:    rdata = 32'hc7d84d1c;
        1331:    rdata = 32'h4d5c8082;
        1332:    rdata = 32'h8082c38c;
        1333:    rdata = 32'hc150c10c;
        1334:    rdata = 32'h010115b7;
        1335:    rdata = 32'h40000613;
        1336:    rdata = 32'ha4890521;
        1337:    rdata = 32'hc5934118;
        1338:    rdata = 32'hf7930015;
        1339:    rdata = 32'h430c0015;
        1340:    rdata = 32'h8ddd99f9;
        1341:    rdata = 32'h8082c30c;
        1342:    rdata = 32'h431c4118;
        1343:    rdata = 32'h0027e793;
        1344:    rdata = 32'h8082c31c;
        1345:    rdata = 32'h4388415c;
        1346:    rdata = 32'h80828905;
        1347:    rdata = 32'hdc227139;
        1348:    rdata = 32'h44334411;
        1349:    rdata = 32'h41180286;
        1350:    rdata = 32'hd84ada26;
        1351:    rdata = 32'hd452d64e;
        1352:    rdata = 32'hce5ed256;
        1353:    rdata = 32'hde06cc62;
        1354:    rdata = 32'h431cd05a;
        1355:    rdata = 32'h89ae84aa;
        1356:    rdata = 32'h89329bf9;
        1357:    rdata = 32'h4a01c31c;
        1358:    rdata = 32'h4c114a81;
        1359:    rdata = 32'h00850b93;
        1360:    rdata = 32'h028ad963;
        1361:    rdata = 32'h86334781;
        1362:    rdata = 32'h06b30149;
        1363:    rdata = 32'hc68300f6;
        1364:    rdata = 32'h00780006;
        1365:    rdata = 32'h0023973e;
        1366:    rdata = 32'h078500d7;
        1367:    rdata = 32'hff8797e3;
        1368:    rdata = 32'h85d24b32;
        1369:    rdata = 32'h22d1855e;
        1370:    rdata = 32'h01652023;
        1371:    rdata = 32'h0a110a85;
        1372:    rdata = 32'h4581bfc1;
        1373:    rdata = 32'h0ab45433;
        1374:    rdata = 32'h00241593;
        1375:    rdata = 32'h40b90533;
        1376:    rdata = 32'h02b90a63;
        1377:    rdata = 32'h468d4781;
        1378:    rdata = 32'hd7634701;
        1379:    rdata = 32'h873300a7;
        1380:    rdata = 32'h974e00f5;
        1381:    rdata = 32'h00074703;
        1382:    rdata = 32'h963e0070;
        1383:    rdata = 32'h00e60023;
        1384:    rdata = 32'h93e30785;
        1385:    rdata = 32'h07a3fed7;
        1386:    rdata = 32'h44320001;
        1387:    rdata = 32'h00848513;
        1388:    rdata = 32'hc1002aad;
        1389:    rdata = 32'h431c4098;
        1390:    rdata = 32'h0017e793;
        1391:    rdata = 32'h50f2c31c;
        1392:    rdata = 32'h54d25462;
        1393:    rdata = 32'h59b25942;
        1394:    rdata = 32'h5a925a22;
        1395:    rdata = 32'h4bf25b02;
        1396:    rdata = 32'h61214c62;
        1397:    rdata = 32'h06138082;
        1398:    rdata = 32'he5910670;
        1399:    rdata = 32'h00000597;
        1400:    rdata = 32'h43058593;
        1401:    rdata = 32'h0597b725;
        1402:    rdata = 32'h85930000;
        1403:    rdata = 32'hbfdd48e5;
        1404:    rdata = 32'h05974625;
        1405:    rdata = 32'h85930000;
        1406:    rdata = 32'hbf094ea5;
        1407:    rdata = 32'h05974625;
        1408:    rdata = 32'h85930000;
        1409:    rdata = 32'hb7194ea5;
        1410:    rdata = 32'h00458793;
        1411:    rdata = 32'hc15cc10c;
        1412:    rdata = 32'h00858793;
        1413:    rdata = 32'hc51c05b1;
        1414:    rdata = 32'h8082c54c;
        1415:    rdata = 32'h431c4118;
        1416:    rdata = 32'h0017e793;
        1417:    rdata = 32'h8082c31c;
        1418:    rdata = 32'h431c4118;
        1419:    rdata = 32'hc31c9bf9;
        1420:    rdata = 32'h41588082;
        1421:    rdata = 32'h9bf9431c;
        1422:    rdata = 32'h8082c31c;
        1423:    rdata = 32'h00458793;
        1424:    rdata = 32'h8793c15c;
        1425:    rdata = 32'hc51c0085;
        1426:    rdata = 32'h00c58793;
        1427:    rdata = 32'h8793c55c;
        1428:    rdata = 32'hc91c0105;
        1429:    rdata = 32'hc10c47b1;
        1430:    rdata = 32'h00f58823;
        1431:    rdata = 32'he793419c;
        1432:    rdata = 32'hc19c0017;
        1433:    rdata = 32'h415c8082;
        1434:    rdata = 32'h8b85439c;
        1435:    rdata = 32'h455cdfed;
        1436:    rdata = 32'h0007c503;
        1437:    rdata = 32'h0ff57513;
        1438:    rdata = 32'h11018082;
        1439:    rdata = 32'hca26cc22;
        1440:    rdata = 32'hc64ec84a;
        1441:    rdata = 32'hc05ac256;
        1442:    rdata = 32'hc452ce06;
        1443:    rdata = 32'h892e84aa;
        1444:    rdata = 32'h440189b2;
        1445:    rdata = 32'h4b214aa9;
        1446:    rdata = 32'h03345f63;
        1447:    rdata = 32'h0a338526;
        1448:    rdata = 32'h37d10089;
        1449:    rdata = 32'h00aa0023;
        1450:    rdata = 32'h01551f63;
        1451:    rdata = 32'h000a0023;
        1452:    rdata = 32'h40f24501;
        1453:    rdata = 32'h44d24462;
        1454:    rdata = 32'h49b24942;
        1455:    rdata = 32'h4a924a22;
        1456:    rdata = 32'h61054b02;
        1457:    rdata = 32'h14638082;
        1458:    rdata = 32'hc4010165;
        1459:    rdata = 32'h04051479;
        1460:    rdata = 32'h547db7e1;
        1461:    rdata = 32'h4505bfed;
        1462:    rdata = 32'h451cbfe9;
        1463:    rdata = 32'h00b78023;
        1464:    rdata = 32'h439c415c;
        1465:    rdata = 32'h4817d793;
        1466:    rdata = 32'h8082ffe5;
        1467:    rdata = 32'hc4221141;
        1468:    rdata = 32'hc606c226;
        1469:    rdata = 32'h842e84aa;
        1470:    rdata = 32'h00044583;
        1471:    rdata = 32'h8526c589;
        1472:    rdata = 32'h3fe10405;
        1473:    rdata = 32'h40b2bfd5;
        1474:    rdata = 32'h44924422;
        1475:    rdata = 32'h80820141;
        1476:    rdata = 32'h4388415c;
        1477:    rdata = 32'h80828905;
        1478:    rdata = 32'hc503455c;
        1479:    rdata = 32'h75130007;
        1480:    rdata = 32'h80820ff5;
        1481:    rdata = 32'hc150c10c;
        1482:    rdata = 32'h41088082;
        1483:    rdata = 32'h952e99f1;
        1484:    rdata = 32'h41488082;
        1485:    rdata = 32'h00008082;
        1486:    rdata = 32'h00a5c7b3;
        1487:    rdata = 32'h0037f793;
        1488:    rdata = 32'h00c508b3;
        1489:    rdata = 32'h06079263;
        1490:    rdata = 32'h00300793;
        1491:    rdata = 32'h04c7fe63;
        1492:    rdata = 32'h00357793;
        1493:    rdata = 32'h00050713;
        1494:    rdata = 32'h06079863;
        1495:    rdata = 32'hffc8f613;
        1496:    rdata = 32'hfe060793;
        1497:    rdata = 32'h08f76c63;
        1498:    rdata = 32'h02c77c63;
        1499:    rdata = 32'h00058693;
        1500:    rdata = 32'h00070793;
        1501:    rdata = 32'h0006a803;
        1502:    rdata = 32'h00478793;
        1503:    rdata = 32'h00468693;
        1504:    rdata = 32'hff07ae23;
        1505:    rdata = 32'hfec7e8e3;
        1506:    rdata = 32'hfff60793;
        1507:    rdata = 32'h40e787b3;
        1508:    rdata = 32'hffc7f793;
        1509:    rdata = 32'h00478793;
        1510:    rdata = 32'h00f70733;
        1511:    rdata = 32'h00f585b3;
        1512:    rdata = 32'h01176863;
        1513:    rdata = 32'h00008067;
        1514:    rdata = 32'h00050713;
        1515:    rdata = 32'hff157ce3;
        1516:    rdata = 32'h0005c783;
        1517:    rdata = 32'h00170713;
        1518:    rdata = 32'h00158593;
        1519:    rdata = 32'hfef70fa3;
        1520:    rdata = 32'hff1768e3;
        1521:    rdata = 32'h00008067;
        1522:    rdata = 32'h0005c683;
        1523:    rdata = 32'h00170713;
        1524:    rdata = 32'h00377793;
        1525:    rdata = 32'hfed70fa3;
        1526:    rdata = 32'h00158593;
        1527:    rdata = 32'hf80780e3;
        1528:    rdata = 32'h0005c683;
        1529:    rdata = 32'h00170713;
        1530:    rdata = 32'h00377793;
        1531:    rdata = 32'hfed70fa3;
        1532:    rdata = 32'h00158593;
        1533:    rdata = 32'hfc079ae3;
        1534:    rdata = 32'hf65ff06f;
        1535:    rdata = 32'h0045a683;
        1536:    rdata = 32'h0005a283;
        1537:    rdata = 32'h0085af83;
        1538:    rdata = 32'h00c5af03;
        1539:    rdata = 32'h0105ae83;
        1540:    rdata = 32'h0145ae03;
        1541:    rdata = 32'h0185a303;
        1542:    rdata = 32'h01c5a803;
        1543:    rdata = 32'h00d72223;
        1544:    rdata = 32'h0205a683;
        1545:    rdata = 32'h00572023;
        1546:    rdata = 32'h01f72423;
        1547:    rdata = 32'h01e72623;
        1548:    rdata = 32'h01d72823;
        1549:    rdata = 32'h01c72a23;
        1550:    rdata = 32'h00672c23;
        1551:    rdata = 32'h01072e23;
        1552:    rdata = 32'h02d72023;
        1553:    rdata = 32'h02470713;
        1554:    rdata = 32'h02458593;
        1555:    rdata = 32'hfaf768e3;
        1556:    rdata = 32'hf19ff06f;
        1557:    rdata = 32'h00f00313;
        1558:    rdata = 32'h00050713;
        1559:    rdata = 32'h02c37e63;
        1560:    rdata = 32'h00f77793;
        1561:    rdata = 32'h0a079063;
        1562:    rdata = 32'h08059263;
        1563:    rdata = 32'hff067693;
        1564:    rdata = 32'h00f67613;
        1565:    rdata = 32'h00e686b3;
        1566:    rdata = 32'h00b72023;
        1567:    rdata = 32'h00b72223;
        1568:    rdata = 32'h00b72423;
        1569:    rdata = 32'h00b72623;
        1570:    rdata = 32'h01070713;
        1571:    rdata = 32'hfed766e3;
        1572:    rdata = 32'h00061463;
        1573:    rdata = 32'h00008067;
        1574:    rdata = 32'h40c306b3;
        1575:    rdata = 32'h00269693;
        1576:    rdata = 32'h00000297;
        1577:    rdata = 32'h005686b3;
        1578:    rdata = 32'h00c68067;
        1579:    rdata = 32'h00b70723;
        1580:    rdata = 32'h00b706a3;
        1581:    rdata = 32'h00b70623;
        1582:    rdata = 32'h00b705a3;
        1583:    rdata = 32'h00b70523;
        1584:    rdata = 32'h00b704a3;
        1585:    rdata = 32'h00b70423;
        1586:    rdata = 32'h00b703a3;
        1587:    rdata = 32'h00b70323;
        1588:    rdata = 32'h00b702a3;
        1589:    rdata = 32'h00b70223;
        1590:    rdata = 32'h00b701a3;
        1591:    rdata = 32'h00b70123;
        1592:    rdata = 32'h00b700a3;
        1593:    rdata = 32'h00b70023;
        1594:    rdata = 32'h00008067;
        1595:    rdata = 32'h0ff5f593;
        1596:    rdata = 32'h00859693;
        1597:    rdata = 32'h00d5e5b3;
        1598:    rdata = 32'h01059693;
        1599:    rdata = 32'h00d5e5b3;
        1600:    rdata = 32'hf6dff06f;
        1601:    rdata = 32'h00279693;
        1602:    rdata = 32'h00000297;
        1603:    rdata = 32'h005686b3;
        1604:    rdata = 32'h00008293;
        1605:    rdata = 32'hfa0680e7;
        1606:    rdata = 32'h00028093;
        1607:    rdata = 32'hff078793;
        1608:    rdata = 32'h40f70733;
        1609:    rdata = 32'h00f60633;
        1610:    rdata = 32'hf6c378e3;
        1611:    rdata = 32'hf3dff06f;
        1612:    rdata = 32'h05971101;
        1613:    rdata = 32'h85930000;
        1614:    rdata = 32'he51766a5;
        1615:    rdata = 32'h0513000e;
        1616:    rdata = 32'hce0674e5;
        1617:    rdata = 32'h80dff0ef;
        1618:    rdata = 32'he0ef0068;
        1619:    rdata = 32'h40f2cf9f;
        1620:    rdata = 32'h61054501;
        1621:    rdata = 32'h05b78082;
        1622:    rdata = 32'he5170100;
        1623:    rdata = 32'h0513000e;
        1624:    rdata = 32'hf06f6b25;
        1625:    rdata = 32'h05b79e3f;
        1626:    rdata = 32'he5170101;
        1627:    rdata = 32'h0513000e;
        1628:    rdata = 32'hf06f6c65;
        1629:    rdata = 32'h37b7ab7f;
        1630:    rdata = 32'he7170100;
        1631:    rdata = 32'h0713000e;
        1632:    rdata = 32'h86936e67;
        1633:    rdata = 32'hc31c0047;
        1634:    rdata = 32'h8693c354;
        1635:    rdata = 32'h07b10087;
        1636:    rdata = 32'hc75cc714;
        1637:    rdata = 32'h25b78082;
        1638:    rdata = 32'he5170100;
        1639:    rdata = 32'h0513000e;
        1640:    rdata = 32'hb9696d65;
        1641:    rdata = 32'h000ee797;
        1642:    rdata = 32'h6e878793;
        1643:    rdata = 32'hc3986741;
        1644:    rdata = 32'hc3d86711;
        1645:    rdata = 32'h00008082;
        1646:    rdata = 32'h00000000;
        1647:    rdata = 32'h00000000;
        1648:    rdata = 32'h00000000;
        1649:    rdata = 32'h00000000;
        1650:    rdata = 32'h00011956;
        1651:    rdata = 32'h00011966;
        1652:    rdata = 32'h00011976;
        1653:    rdata = 32'h00011996;
        1654:    rdata = 32'h000119a4;
        1655:    rdata = 32'hffffecdc;
        1656:    rdata = 32'hffffece2;
        1657:    rdata = 32'hffffece8;
        1658:    rdata = 32'hffffecee;
        1659:    rdata = 32'hffffecfc;
        1660:    rdata = 32'hffffed04;
        1661:    rdata = 32'hffffed0c;
        1662:    rdata = 32'hffffed14;
        1663:    rdata = 32'hffffed1c;
        1664:    rdata = 32'hffffed24;
        1665:    rdata = 32'hffffed2a;
        1666:    rdata = 32'hffffed30;
        1667:    rdata = 32'h0002c000;
        1668:    rdata = 32'h0003c000;
        1669:    rdata = 32'hc00002c0;
        1670:    rdata = 32'h02c00003;
        1671:    rdata = 32'h0003c000;
        1672:    rdata = 32'hc00002c0;
        1673:    rdata = 32'h02c00003;
        1674:    rdata = 32'h0003c000;
        1675:    rdata = 32'hc00002c0;
        1676:    rdata = 32'h02c00003;
        1677:    rdata = 32'h0003c000;
        1678:    rdata = 32'hc00002c0;
        1679:    rdata = 32'h02c00003;
        1680:    rdata = 32'h0003c000;
        1681:    rdata = 32'hc00002c0;
        1682:    rdata = 32'h02c00003;
        1683:    rdata = 32'h0003c000;
        1684:    rdata = 32'hc00002c0;
        1685:    rdata = 32'h02c00003;
        1686:    rdata = 32'h0003c000;
        1687:    rdata = 32'hc00002c0;
        1688:    rdata = 32'h02c00003;
        1689:    rdata = 32'h0003c000;
        1690:    rdata = 32'hc00002c0;
        1691:    rdata = 32'h02c00003;
        1692:    rdata = 32'h00042000;
        1693:    rdata = 32'h0002c000;
        1694:    rdata = 32'h0005c000;
        1695:    rdata = 32'hc00004c0;
        1696:    rdata = 32'h04c00005;
        1697:    rdata = 32'h0005c000;
        1698:    rdata = 32'hc00004c0;
        1699:    rdata = 32'h04c00005;
        1700:    rdata = 32'h0005c000;
        1701:    rdata = 32'hc00004c0;
        1702:    rdata = 32'h04c00005;
        1703:    rdata = 32'h0005c000;
        1704:    rdata = 32'hc00004c0;
        1705:    rdata = 32'h04c00005;
        1706:    rdata = 32'h0005c000;
        1707:    rdata = 32'hc00004c0;
        1708:    rdata = 32'h04c00005;
        1709:    rdata = 32'h0005c000;
        1710:    rdata = 32'hc00004c0;
        1711:    rdata = 32'h04c00005;
        1712:    rdata = 32'h0005c000;
        1713:    rdata = 32'hc00004c0;
        1714:    rdata = 32'h04c00005;
        1715:    rdata = 32'h0005c000;
        1716:    rdata = 32'hc00004c0;
        1717:    rdata = 32'h04c00005;
        1718:    rdata = 32'h00042000;
        1719:    rdata = 32'h0020c000;
        1720:    rdata = 32'h200000c0;
        1721:    rdata = 32'h00000000;
        1722:    rdata = 32'h0008c000;
        1723:    rdata = 32'h200000c0;
        1724:    rdata = 32'h00000000;
        1725:    rdata = 32'h72616568;
        1726:    rdata = 32'h61656274;
        1727:    rdata = 32'h00000a74;
        1728:    rdata = 32'h706c6568;
        1729:    rdata = 32'h20202020;
        1730:    rdata = 32'h20202020;
        1731:    rdata = 32'h20202020;
        1732:    rdata = 32'h20202020;
        1733:    rdata = 32'h20202020;
        1734:    rdata = 32'h20202020;
        1735:    rdata = 32'h20202020;
        1736:    rdata = 32'h202d2020;
        1737:    rdata = 32'h6e697270;
        1738:    rdata = 32'h68742074;
        1739:    rdata = 32'h6d207369;
        1740:    rdata = 32'h61737365;
        1741:    rdata = 32'h720a6567;
        1742:    rdata = 32'h74657365;
        1743:    rdata = 32'h20202020;
        1744:    rdata = 32'h20202020;
        1745:    rdata = 32'h20202020;
        1746:    rdata = 32'h20202020;
        1747:    rdata = 32'h20202020;
        1748:    rdata = 32'h20202020;
        1749:    rdata = 32'h20202020;
        1750:    rdata = 32'h72202d20;
        1751:    rdata = 32'h74657365;
        1752:    rdata = 32'h636f7320;
        1753:    rdata = 32'h6e69700a;
        1754:    rdata = 32'h20202067;
        1755:    rdata = 32'h20202020;
        1756:    rdata = 32'h20202020;
        1757:    rdata = 32'h20202020;
        1758:    rdata = 32'h20202020;
        1759:    rdata = 32'h20202020;
        1760:    rdata = 32'h20202020;
        1761:    rdata = 32'h2d202020;
        1762:    rdata = 32'h6e657320;
        1763:    rdata = 32'h70222064;
        1764:    rdata = 32'h22676e69;
        1765:    rdata = 32'h206f7420;
        1766:    rdata = 32'h20656874;
        1767:    rdata = 32'h74736f68;
        1768:    rdata = 32'h7465730a;
        1769:    rdata = 32'h6970675f;
        1770:    rdata = 32'h69645f6f;
        1771:    rdata = 32'h74636572;
        1772:    rdata = 32'h206e6f69;
        1773:    rdata = 32'h6e69703c;
        1774:    rdata = 32'h695b203e;
        1775:    rdata = 32'h756f7c6e;
        1776:    rdata = 32'h2d205d74;
        1777:    rdata = 32'h74657320;
        1778:    rdata = 32'h69706720;
        1779:    rdata = 32'h6970206f;
        1780:    rdata = 32'h6964206e;
        1781:    rdata = 32'h74636572;
        1782:    rdata = 32'h0a6e6f69;
        1783:    rdata = 32'h5f746567;
        1784:    rdata = 32'h6f697067;
        1785:    rdata = 32'h7269645f;
        1786:    rdata = 32'h69746365;
        1787:    rdata = 32'h3c206e6f;
        1788:    rdata = 32'h3e6e6970;
        1789:    rdata = 32'h20202020;
        1790:    rdata = 32'h20202020;
        1791:    rdata = 32'h202d2020;
        1792:    rdata = 32'h20746567;
        1793:    rdata = 32'h6f697067;
        1794:    rdata = 32'h6e697020;
        1795:    rdata = 32'h72696420;
        1796:    rdata = 32'h69746365;
        1797:    rdata = 32'h730a6e6f;
        1798:    rdata = 32'h675f7465;
        1799:    rdata = 32'h206f6970;
        1800:    rdata = 32'h6e69703c;
        1801:    rdata = 32'h763c203e;
        1802:    rdata = 32'h65756c61;
        1803:    rdata = 32'h2020203e;
        1804:    rdata = 32'h20202020;
        1805:    rdata = 32'h20202020;
        1806:    rdata = 32'h73202d20;
        1807:    rdata = 32'h67207465;
        1808:    rdata = 32'h206f6970;
        1809:    rdata = 32'h0a6e6970;
        1810:    rdata = 32'h5f746567;
        1811:    rdata = 32'h6f697067;
        1812:    rdata = 32'h69703c20;
        1813:    rdata = 32'h20203e6e;
        1814:    rdata = 32'h20202020;
        1815:    rdata = 32'h20202020;
        1816:    rdata = 32'h20202020;
        1817:    rdata = 32'h20202020;
        1818:    rdata = 32'h202d2020;
        1819:    rdata = 32'h20746567;
        1820:    rdata = 32'h6f697067;
        1821:    rdata = 32'h6e697020;
        1822:    rdata = 32'h7465730a;
        1823:    rdata = 32'h6165685f;
        1824:    rdata = 32'h65627472;
        1825:    rdata = 32'h3c207461;
        1826:    rdata = 32'h69726570;
        1827:    rdata = 32'h5b20646f;
        1828:    rdata = 32'h3e5d736d;
        1829:    rdata = 32'h20202020;
        1830:    rdata = 32'h2d202020;
        1831:    rdata = 32'h74657320;
        1832:    rdata = 32'h61656820;
        1833:    rdata = 32'h65627472;
        1834:    rdata = 32'h630a7461;
        1835:    rdata = 32'h75636c61;
        1836:    rdata = 32'h6574616c;
        1837:    rdata = 32'h72613c20;
        1838:    rdata = 32'h203e3167;
        1839:    rdata = 32'h2d7c2b5b;
        1840:    rdata = 32'h2f7c2a7c;
        1841:    rdata = 32'h613c205d;
        1842:    rdata = 32'h3e326772;
        1843:    rdata = 32'h70202d20;
        1844:    rdata = 32'h6f667265;
        1845:    rdata = 32'h63206d72;
        1846:    rdata = 32'h75636c61;
        1847:    rdata = 32'h6974616c;
        1848:    rdata = 32'h720a6e6f;
        1849:    rdata = 32'h5f646165;
        1850:    rdata = 32'h7274616d;
        1851:    rdata = 32'h20207869;
        1852:    rdata = 32'h20202020;
        1853:    rdata = 32'h20202020;
        1854:    rdata = 32'h20202020;
        1855:    rdata = 32'h20202020;
        1856:    rdata = 32'h20202020;
        1857:    rdata = 32'h72202d20;
        1858:    rdata = 32'h20646165;
        1859:    rdata = 32'h7274616d;
        1860:    rdata = 32'h630a7869;
        1861:    rdata = 32'h62696c61;
        1862:    rdata = 32'h65746172;
        1863:    rdata = 32'h74616d5f;
        1864:    rdata = 32'h20786972;
        1865:    rdata = 32'h20202020;
        1866:    rdata = 32'h20202020;
        1867:    rdata = 32'h20202020;
        1868:    rdata = 32'h20202020;
        1869:    rdata = 32'h63202d20;
        1870:    rdata = 32'h62696c61;
        1871:    rdata = 32'h65746172;
        1872:    rdata = 32'h78697020;
        1873:    rdata = 32'h20736c65;
        1874:    rdata = 32'h7366666f;
        1875:    rdata = 32'h0a737465;
        1876:    rdata = 32'h00000000;
        1877:    rdata = 32'h6f727265;
        1878:    rdata = 32'h6f203a72;
        1879:    rdata = 32'h61726570;
        1880:    rdata = 32'h6e6f6974;
        1881:    rdata = 32'h746f6e20;
        1882:    rdata = 32'h70757320;
        1883:    rdata = 32'h74726f70;
        1884:    rdata = 32'h000a6465;
        1885:    rdata = 32'h676e6970;
        1886:    rdata = 32'h0000000a;
        1887:    rdata = 32'h6f727265;
        1888:    rdata = 32'h6d203a72;
        1889:    rdata = 32'h69737369;
        1890:    rdata = 32'h6120676e;
        1891:    rdata = 32'h6d756772;
        1892:    rdata = 32'h28746e65;
        1893:    rdata = 32'h000a2973;
        1894:    rdata = 32'h6f727265;
        1895:    rdata = 32'h69203a72;
        1896:    rdata = 32'h6c61766e;
        1897:    rdata = 32'h61206469;
        1898:    rdata = 32'h6d756772;
        1899:    rdata = 32'h28746e65;
        1900:    rdata = 32'h74202973;
        1901:    rdata = 32'h28657079;
        1902:    rdata = 32'h000a2973;
        1903:    rdata = 32'h00006e69;
        1904:    rdata = 32'h0074756f;
        1905:    rdata = 32'h6f727265;
        1906:    rdata = 32'h69203a72;
        1907:    rdata = 32'h6c61766e;
        1908:    rdata = 32'h64206469;
        1909:    rdata = 32'h63657269;
        1910:    rdata = 32'h6e6f6974;
        1911:    rdata = 32'h0000000a;
        1912:    rdata = 32'h6f727265;
        1913:    rdata = 32'h6d203a72;
        1914:    rdata = 32'h69737369;
        1915:    rdata = 32'h6120676e;
        1916:    rdata = 32'h6d756772;
        1917:    rdata = 32'h0a746e65;
        1918:    rdata = 32'h00000000;
        1919:    rdata = 32'h6f727265;
        1920:    rdata = 32'h69203a72;
        1921:    rdata = 32'h6c61766e;
        1922:    rdata = 32'h61206469;
        1923:    rdata = 32'h6d756772;
        1924:    rdata = 32'h20746e65;
        1925:    rdata = 32'h65707974;
        1926:    rdata = 32'h0000000a;
        1927:    rdata = 32'h6f727265;
        1928:    rdata = 32'h64203a72;
        1929:    rdata = 32'h73697669;
        1930:    rdata = 32'h206e6f69;
        1931:    rdata = 32'h7a207962;
        1932:    rdata = 32'h0a6f7265;
        1933:    rdata = 32'h00000000;
        1934:    rdata = 32'h6f727265;
        1935:    rdata = 32'h75203a72;
        1936:    rdata = 32'h6365726e;
        1937:    rdata = 32'h696e676f;
        1938:    rdata = 32'h2064657a;
        1939:    rdata = 32'h7265706f;
        1940:    rdata = 32'h6f697461;
        1941:    rdata = 32'h00000a6e;
        1942:    rdata = 32'h64616572;
        1943:    rdata = 32'h5f74756f;
        1944:    rdata = 32'h656d6974;
        1945:    rdata = 32'h00000000;
        1946:    rdata = 32'h7366666f;
        1947:    rdata = 32'h63207465;
        1948:    rdata = 32'h62696c61;
        1949:    rdata = 32'h69746172;
        1950:    rdata = 32'h64206e6f;
        1951:    rdata = 32'h0a656e6f;
        1952:    rdata = 32'h00000000;
        1953:    rdata = 32'h696c6163;
        1954:    rdata = 32'h74617262;
        1955:    rdata = 32'h5f6e6f69;
        1956:    rdata = 32'h656d6974;
        1957:    rdata = 32'h00000000;
        1958:    rdata = 32'h0000203e;
        1959:    rdata = 32'h6f727265;
        1960:    rdata = 32'h75203a72;
        1961:    rdata = 32'h6365726e;
        1962:    rdata = 32'h696e676f;
        1963:    rdata = 32'h2064657a;
        1964:    rdata = 32'h6d6d6f63;
        1965:    rdata = 32'h3a646e61;
        1966:    rdata = 32'h00002220;
        1967:    rdata = 32'h65202e22;
        1968:    rdata = 32'h75636578;
        1969:    rdata = 32'h22206574;
        1970:    rdata = 32'h706c6568;
        1971:    rdata = 32'h6f742022;
        1972:    rdata = 32'h74656720;
        1973:    rdata = 32'h70757320;
        1974:    rdata = 32'h74726f70;
        1975:    rdata = 32'h63206465;
        1976:    rdata = 32'h616d6d6f;
        1977:    rdata = 32'h2073646e;
        1978:    rdata = 32'h7473696c;
        1979:    rdata = 32'h0000000a;
        1980:    rdata = 32'h6f727265;
        1981:    rdata = 32'h63203a72;
        1982:    rdata = 32'h616d6d6f;
        1983:    rdata = 32'h6620646e;
        1984:    rdata = 32'h656c6961;
        1985:    rdata = 32'h00000a64;
        1986:    rdata = 32'h706c6568;
        1987:    rdata = 32'h00000000;
        1988:    rdata = 32'h65736572;
        1989:    rdata = 32'h00000074;
        1990:    rdata = 32'h676e6970;
        1991:    rdata = 32'h00000000;
        1992:    rdata = 32'h5f746573;
        1993:    rdata = 32'h6f697067;
        1994:    rdata = 32'h7269645f;
        1995:    rdata = 32'h69746365;
        1996:    rdata = 32'h00006e6f;
        1997:    rdata = 32'h5f746567;
        1998:    rdata = 32'h6f697067;
        1999:    rdata = 32'h7269645f;
        2000:    rdata = 32'h69746365;
        2001:    rdata = 32'h00006e6f;
        2002:    rdata = 32'h5f746573;
        2003:    rdata = 32'h6f697067;
        2004:    rdata = 32'h00000000;
        2005:    rdata = 32'h5f746567;
        2006:    rdata = 32'h6f697067;
        2007:    rdata = 32'h00000000;
        2008:    rdata = 32'h5f746573;
        2009:    rdata = 32'h72616568;
        2010:    rdata = 32'h61656274;
        2011:    rdata = 32'h00000074;
        2012:    rdata = 32'h636c6163;
        2013:    rdata = 32'h74616c75;
        2014:    rdata = 32'h00000065;
        2015:    rdata = 32'h64616572;
        2016:    rdata = 32'h74616d5f;
        2017:    rdata = 32'h00786972;
        2018:    rdata = 32'h696c6163;
        2019:    rdata = 32'h74617262;
        2020:    rdata = 32'h616d5f65;
        2021:    rdata = 32'h78697274;
        2022:    rdata = 32'h00000000;
        2023:    rdata = 32'h6d6d6f63;
        2024:    rdata = 32'h5f646e61;
        2025:    rdata = 32'h65746e69;
        2026:    rdata = 32'h65727072;
        2027:    rdata = 32'h20726574;
        2028:    rdata = 32'h72617473;
        2029:    rdata = 32'h0a646574;
        2030:    rdata = 32'h00000000;
        2031:    rdata = 32'h0000203a;
        2032:    rdata = 32'h00002820;
        2033:    rdata = 32'h00203a29;
        2034:    rdata = 32'h6f636e69;
        2035:    rdata = 32'h63657272;
        2036:    rdata = 32'h61762074;
        2037:    rdata = 32'h2e65756c;
        2038:    rdata = 32'h79727420;
        2039:    rdata = 32'h61676120;
        2040:    rdata = 32'h000a6e69;
        default: rdata = 32'h00000000;
    endcase
end
endmodule
