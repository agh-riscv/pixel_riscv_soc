/**
 * Copyright (C) 2020  AGH University of Science and Technology
 *
 * This program is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with this program.  If not, see <https://www.gnu.org/licenses/>.
 */

module boot_mem (
    output logic [31:0] rdata,
    input logic [31:0] addr
);

/**
 * Module internal logic
 */

always_comb begin
    case (addr[13:2])
           0:    rdata = 32'h08c0006f;
           1:    rdata = 32'h0880006f;
           2:    rdata = 32'h0840006f;
           3:    rdata = 32'h0800006f;
           4:    rdata = 32'h07c0006f;
           5:    rdata = 32'h0780006f;
           6:    rdata = 32'h0740006f;
           7:    rdata = 32'h0700006f;
           8:    rdata = 32'h06c0006f;
           9:    rdata = 32'h0680006f;
          10:    rdata = 32'h0640006f;
          11:    rdata = 32'h0600006f;
          12:    rdata = 32'h05c0006f;
          13:    rdata = 32'h0580006f;
          14:    rdata = 32'h0540006f;
          15:    rdata = 32'h0500006f;
          16:    rdata = 32'h04c0006f;
          17:    rdata = 32'h0480006f;
          18:    rdata = 32'h0440006f;
          19:    rdata = 32'h0400006f;
          20:    rdata = 32'h03c0006f;
          21:    rdata = 32'h0380006f;
          22:    rdata = 32'h0340006f;
          23:    rdata = 32'h0300006f;
          24:    rdata = 32'h02c0006f;
          25:    rdata = 32'h0280006f;
          26:    rdata = 32'h0240006f;
          27:    rdata = 32'h0200006f;
          28:    rdata = 32'h01c0006f;
          29:    rdata = 32'h0180006f;
          30:    rdata = 32'h0140006f;
          31:    rdata = 32'h0100006f;
          32:    rdata = 32'h0100006f;
          33:    rdata = 32'h0080006f;
          34:    rdata = 32'h0040006f;
          35:    rdata = 32'h0000006f;
          36:    rdata = 32'h00000093;
          37:    rdata = 32'h00000113;
          38:    rdata = 32'h00000193;
          39:    rdata = 32'h00000213;
          40:    rdata = 32'h00000293;
          41:    rdata = 32'h00000313;
          42:    rdata = 32'h00000393;
          43:    rdata = 32'h00000413;
          44:    rdata = 32'h00000493;
          45:    rdata = 32'h00000513;
          46:    rdata = 32'h00000593;
          47:    rdata = 32'h00000613;
          48:    rdata = 32'h00000693;
          49:    rdata = 32'h00000713;
          50:    rdata = 32'h00000793;
          51:    rdata = 32'h00000813;
          52:    rdata = 32'h00000893;
          53:    rdata = 32'h00000913;
          54:    rdata = 32'h00000993;
          55:    rdata = 32'h00000a13;
          56:    rdata = 32'h00000a93;
          57:    rdata = 32'h00000b13;
          58:    rdata = 32'h00000b93;
          59:    rdata = 32'h00000c13;
          60:    rdata = 32'h00000c93;
          61:    rdata = 32'h00000d13;
          62:    rdata = 32'h00000d93;
          63:    rdata = 32'h00000e13;
          64:    rdata = 32'h00000e93;
          65:    rdata = 32'h00000f13;
          66:    rdata = 32'h00000f93;
          67:    rdata = 32'h00104117;
          68:    rdata = 32'hef410113;
          69:    rdata = 32'h00100297;
          70:    rdata = 32'heec28293;
          71:    rdata = 32'h00100317;
          72:    rdata = 32'hf3430313;
          73:    rdata = 32'h0062d863;
          74:    rdata = 32'h0002a023;
          75:    rdata = 32'h00428293;
          76:    rdata = 32'hfe535ce3;
          77:    rdata = 32'h5f000293;
          78:    rdata = 32'h00100317;
          79:    rdata = 32'hec830313;
          80:    rdata = 32'h00100397;
          81:    rdata = 32'hec038393;
          82:    rdata = 32'h00735c63;
          83:    rdata = 32'h0002ae03;
          84:    rdata = 32'h01c32023;
          85:    rdata = 32'h00428293;
          86:    rdata = 32'h00430313;
          87:    rdata = 32'hfe7348e3;
          88:    rdata = 32'h55c00293;
          89:    rdata = 32'h56c00313;
          90:    rdata = 32'h0062da63;
          91:    rdata = 32'h0002a783;
          92:    rdata = 32'h000780e7;
          93:    rdata = 32'h00428293;
          94:    rdata = 32'hfe62cae3;
          95:    rdata = 32'h00000513;
          96:    rdata = 32'h00000593;
          97:    rdata = 32'h2d8000ef;
          98:    rdata = 32'h45857179;
          99:    rdata = 32'h00100517;
         100:    rdata = 32'he9450513;
         101:    rdata = 32'hd422d606;
         102:    rdata = 32'hce4ed04a;
         103:    rdata = 32'hd226cc52;
         104:    rdata = 32'h458d2249;
         105:    rdata = 32'h00100517;
         106:    rdata = 32'he7c50513;
         107:    rdata = 32'h44012a61;
         108:    rdata = 32'h00100917;
         109:    rdata = 32'he9890913;
         110:    rdata = 32'h00100997;
         111:    rdata = 32'he6898993;
         112:    rdata = 32'h854a4a11;
         113:    rdata = 32'h73632065;
         114:    rdata = 32'h448102a4;
         115:    rdata = 32'h2abd854e;
         116:    rdata = 32'h97a6007c;
         117:    rdata = 32'h00a78023;
         118:    rdata = 32'h99e30485;
         119:    rdata = 32'h44b2ff44;
         120:    rdata = 32'h854a85a2;
         121:    rdata = 32'hc1042041;
         122:    rdata = 32'hbfe10411;
         123:    rdata = 32'h542250b2;
         124:    rdata = 32'h59025492;
         125:    rdata = 32'h4a6249f2;
         126:    rdata = 32'h80826145;
         127:    rdata = 32'hd4227179;
         128:    rdata = 32'hce4ed04a;
         129:    rdata = 32'hd606cc52;
         130:    rdata = 32'h4401d226;
         131:    rdata = 32'h00100917;
         132:    rdata = 32'he3c90913;
         133:    rdata = 32'h00100997;
         134:    rdata = 32'he2098993;
         135:    rdata = 32'h854a4a11;
         136:    rdata = 32'h736320b1;
         137:    rdata = 32'h448102a4;
         138:    rdata = 32'h2a41854e;
         139:    rdata = 32'h97a6007c;
         140:    rdata = 32'h00a78023;
         141:    rdata = 32'h99e30485;
         142:    rdata = 32'h44b2ff44;
         143:    rdata = 32'h854a85a2;
         144:    rdata = 32'hc1042015;
         145:    rdata = 32'hbfe10411;
         146:    rdata = 32'h542250b2;
         147:    rdata = 32'h59025492;
         148:    rdata = 32'h4a6249f2;
         149:    rdata = 32'h80826145;
         150:    rdata = 32'hb73de111;
         151:    rdata = 32'hc10cb745;
         152:    rdata = 32'h8082c150;
         153:    rdata = 32'h99f14108;
         154:    rdata = 32'h8082952e;
         155:    rdata = 32'h80824148;
         156:    rdata = 32'h00458793;
         157:    rdata = 32'h8793c15c;
         158:    rdata = 32'hc51c0085;
         159:    rdata = 32'h00c58793;
         160:    rdata = 32'h8793c55c;
         161:    rdata = 32'hc91c0105;
         162:    rdata = 32'h01458793;
         163:    rdata = 32'hc95cc10c;
         164:    rdata = 32'h01858793;
         165:    rdata = 32'hcd1c05f1;
         166:    rdata = 32'h8082cd4c;
         167:    rdata = 32'h4388455c;
         168:    rdata = 32'h97b34785;
         169:    rdata = 32'h8d7d00b7;
         170:    rdata = 32'h00a03533;
         171:    rdata = 32'h451c8082;
         172:    rdata = 32'h8e3d439c;
         173:    rdata = 32'h8e3d8e6d;
         174:    rdata = 32'hc390451c;
         175:    rdata = 32'h47858082;
         176:    rdata = 32'h00b61633;
         177:    rdata = 32'h00b795b3;
         178:    rdata = 32'h1141b7dd;
         179:    rdata = 32'hc226c422;
         180:    rdata = 32'h842ac606;
         181:    rdata = 32'h37d984ae;
         182:    rdata = 32'h00154613;
         183:    rdata = 32'h44228522;
         184:    rdata = 32'h85a640b2;
         185:    rdata = 32'h76134492;
         186:    rdata = 32'h01410ff6;
         187:    rdata = 32'h455cbfc9;
         188:    rdata = 32'h55134388;
         189:    rdata = 32'h80824915;
         190:    rdata = 32'h4388455c;
         191:    rdata = 32'h49055513;
         192:    rdata = 32'h862e8082;
         193:    rdata = 32'hbf6545bd;
         194:    rdata = 32'h00458793;
         195:    rdata = 32'h8793c15c;
         196:    rdata = 32'hc10c0085;
         197:    rdata = 32'h8793c51c;
         198:    rdata = 32'h05c100c5;
         199:    rdata = 32'hc90cc55c;
         200:    rdata = 32'h41188082;
         201:    rdata = 32'h0015f793;
         202:    rdata = 32'h99f9430c;
         203:    rdata = 32'hc30c8ddd;
         204:    rdata = 32'h41188082;
         205:    rdata = 32'h97938985;
         206:    rdata = 32'h430c0015;
         207:    rdata = 32'h8ddd99f5;
         208:    rdata = 32'h8082c30c;
         209:    rdata = 32'h8023491c;
         210:    rdata = 32'h808200b7;
         211:    rdata = 32'h8023451c;
         212:    rdata = 32'h415c0007;
         213:    rdata = 32'h8b85439c;
         214:    rdata = 32'h455cdfed;
         215:    rdata = 32'h0007c503;
         216:    rdata = 32'h0ff57513;
         217:    rdata = 32'h451c8082;
         218:    rdata = 32'h00b78023;
         219:    rdata = 32'h439c415c;
         220:    rdata = 32'h4817d793;
         221:    rdata = 32'h455cffe5;
         222:    rdata = 32'h0007c783;
         223:    rdata = 32'h415c8082;
         224:    rdata = 32'h89054388;
         225:    rdata = 32'h415c8082;
         226:    rdata = 32'h55134388;
         227:    rdata = 32'h80824815;
         228:    rdata = 32'h00458793;
         229:    rdata = 32'h8793c15c;
         230:    rdata = 32'hc51c0085;
         231:    rdata = 32'h00c58793;
         232:    rdata = 32'h8793c55c;
         233:    rdata = 32'hc91c0105;
         234:    rdata = 32'hc10c4799;
         235:    rdata = 32'h00f58823;
         236:    rdata = 32'he793419c;
         237:    rdata = 32'hc19c0017;
         238:    rdata = 32'h415c8082;
         239:    rdata = 32'h8b85439c;
         240:    rdata = 32'h455cdfed;
         241:    rdata = 32'h0007c503;
         242:    rdata = 32'h0ff57513;
         243:    rdata = 32'h11018082;
         244:    rdata = 32'hca26cc22;
         245:    rdata = 32'hc64ec84a;
         246:    rdata = 32'hce06c256;
         247:    rdata = 32'h84aac452;
         248:    rdata = 32'h89b2892e;
         249:    rdata = 32'h4aa94401;
         250:    rdata = 32'h03345863;
         251:    rdata = 32'h0a338526;
         252:    rdata = 32'h37e10089;
         253:    rdata = 32'h00aa0023;
         254:    rdata = 32'h01551e63;
         255:    rdata = 32'h000a0023;
         256:    rdata = 32'h40f24501;
         257:    rdata = 32'h44d24462;
         258:    rdata = 32'h49b24942;
         259:    rdata = 32'h4a924a22;
         260:    rdata = 32'h80826105;
         261:    rdata = 32'hbfc90405;
         262:    rdata = 32'hb7e54505;
         263:    rdata = 32'h8023451c;
         264:    rdata = 32'h415c00b7;
         265:    rdata = 32'hd793439c;
         266:    rdata = 32'hffe54817;
         267:    rdata = 32'h11418082;
         268:    rdata = 32'hc226c422;
         269:    rdata = 32'h84aac606;
         270:    rdata = 32'h4583842e;
         271:    rdata = 32'h85260004;
         272:    rdata = 32'h3fe90405;
         273:    rdata = 32'hfff44783;
         274:    rdata = 32'h40b2fbed;
         275:    rdata = 32'h44924422;
         276:    rdata = 32'h80820141;
         277:    rdata = 32'h4388415c;
         278:    rdata = 32'h80828905;
         279:    rdata = 32'h05971141;
         280:    rdata = 32'h85930000;
         281:    rdata = 32'h051710e5;
         282:    rdata = 32'h05130010;
         283:    rdata = 32'hc606bce5;
         284:    rdata = 32'h3f75c422;
         285:    rdata = 32'h00100517;
         286:    rdata = 32'hb8c50513;
         287:    rdata = 32'h05973d8d;
         288:    rdata = 32'h85930000;
         289:    rdata = 32'he91d1025;
         290:    rdata = 32'h00100517;
         291:    rdata = 32'hb7850513;
         292:    rdata = 32'h842a35a5;
         293:    rdata = 32'h00000597;
         294:    rdata = 32'h10058593;
         295:    rdata = 32'h0597e509;
         296:    rdata = 32'h85930000;
         297:    rdata = 32'h051710e5;
         298:    rdata = 32'h05130010;
         299:    rdata = 32'h3741b8e5;
         300:    rdata = 32'h335d8522;
         301:    rdata = 32'h00000597;
         302:    rdata = 32'h11058593;
         303:    rdata = 32'h00100517;
         304:    rdata = 32'hb7850513;
         305:    rdata = 32'h62c137ad;
         306:    rdata = 32'h305292f3;
         307:    rdata = 32'h00000597;
         308:    rdata = 32'h10c58593;
         309:    rdata = 32'h00100517;
         310:    rdata = 32'hb6050513;
         311:    rdata = 32'h45853f89;
         312:    rdata = 32'h00100517;
         313:    rdata = 32'hb2050513;
         314:    rdata = 32'hf06f3d29;
         315:    rdata = 32'h40b23970;
         316:    rdata = 32'h45014422;
         317:    rdata = 32'h80820141;
         318:    rdata = 32'h00100797;
         319:    rdata = 32'hb5078793;
         320:    rdata = 32'hc3986741;
         321:    rdata = 32'hc3d86711;
         322:    rdata = 32'h05b78082;
         323:    rdata = 32'h05170100;
         324:    rdata = 32'h05130010;
         325:    rdata = 32'hbba9af25;
         326:    rdata = 32'h010017b7;
         327:    rdata = 32'h00100717;
         328:    rdata = 32'hb0470713;
         329:    rdata = 32'h00478693;
         330:    rdata = 32'h8693c354;
         331:    rdata = 32'hc31c0087;
         332:    rdata = 32'h8693c714;
         333:    rdata = 32'h07c100c7;
         334:    rdata = 32'hcb1cc754;
         335:    rdata = 32'h25b78082;
         336:    rdata = 32'h05170100;
         337:    rdata = 32'h05130010;
         338:    rdata = 32'hb599af25;
         339:    rdata = 32'h00000000;
         340:    rdata = 32'h00000000;
         341:    rdata = 32'h00000000;
         342:    rdata = 32'h00000000;
         343:    rdata = 32'h000004f8;
         344:    rdata = 32'h0000050a;
         345:    rdata = 32'h00000518;
         346:    rdata = 32'h0000053e;
         347:    rdata = 32'h746f6f62;
         348:    rdata = 32'h64616f6c;
         349:    rdata = 32'h73207265;
         350:    rdata = 32'h74726174;
         351:    rdata = 32'h000a6465;
         352:    rdata = 32'h65646f63;
         353:    rdata = 32'h64616f6c;
         354:    rdata = 32'h696b7320;
         355:    rdata = 32'h64657070;
         356:    rdata = 32'h0000000a;
         357:    rdata = 32'h65646f63;
         358:    rdata = 32'h64616f6c;
         359:    rdata = 32'h756f7320;
         360:    rdata = 32'h3a656372;
         361:    rdata = 32'h72617520;
         362:    rdata = 32'h00000a74;
         363:    rdata = 32'h65646f63;
         364:    rdata = 32'h64616f6c;
         365:    rdata = 32'h756f7320;
         366:    rdata = 32'h3a656372;
         367:    rdata = 32'h69707320;
         368:    rdata = 32'h0000000a;
         369:    rdata = 32'h65646f63;
         370:    rdata = 32'h64616f6c;
         371:    rdata = 32'h6e696620;
         372:    rdata = 32'h65687369;
         373:    rdata = 32'h00000a64;
         374:    rdata = 32'h746f6f62;
         375:    rdata = 32'h64616f6c;
         376:    rdata = 32'h66207265;
         377:    rdata = 32'h73696e69;
         378:    rdata = 32'h0a646568;
         379:    rdata = 32'h00000000;
        default: rdata = 32'h00000000;
    endcase
end
endmodule
