/**
 * Copyright (C) 2020  AGH University of Science and Technology
 *
 * This program is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with this program.  If not, see <https://www.gnu.org/licenses/>.
 */

module spi_mem (
    output logic [31:0] rdata,
    input logic [31:0] addr
);

/**
 * Module internal logic
 */

always_comb begin
    case (addr[13:2])
           0:    rdata = 32'h08c0006f;
           1:    rdata = 32'h0880006f;
           2:    rdata = 32'h0840006f;
           3:    rdata = 32'h0800006f;
           4:    rdata = 32'h07c0006f;
           5:    rdata = 32'h0780006f;
           6:    rdata = 32'h0740006f;
           7:    rdata = 32'h0700006f;
           8:    rdata = 32'h06c0006f;
           9:    rdata = 32'h0680006f;
          10:    rdata = 32'h0640006f;
          11:    rdata = 32'h0600006f;
          12:    rdata = 32'h05c0006f;
          13:    rdata = 32'h0580006f;
          14:    rdata = 32'h0540006f;
          15:    rdata = 32'h0500006f;
          16:    rdata = 32'h3510006f;
          17:    rdata = 32'h39f0006f;
          18:    rdata = 32'h0440006f;
          19:    rdata = 32'h0400006f;
          20:    rdata = 32'h03c0006f;
          21:    rdata = 32'h0380006f;
          22:    rdata = 32'h0340006f;
          23:    rdata = 32'h0300006f;
          24:    rdata = 32'h02c0006f;
          25:    rdata = 32'h0280006f;
          26:    rdata = 32'h0240006f;
          27:    rdata = 32'h0200006f;
          28:    rdata = 32'h01c0006f;
          29:    rdata = 32'h0180006f;
          30:    rdata = 32'h0140006f;
          31:    rdata = 32'h0100006f;
          32:    rdata = 32'h0100006f;
          33:    rdata = 32'h0080006f;
          34:    rdata = 32'h0040006f;
          35:    rdata = 32'h0000006f;
          36:    rdata = 32'h00000093;
          37:    rdata = 32'h00000113;
          38:    rdata = 32'h00000193;
          39:    rdata = 32'h00000213;
          40:    rdata = 32'h00000293;
          41:    rdata = 32'h00000313;
          42:    rdata = 32'h00000393;
          43:    rdata = 32'h00000413;
          44:    rdata = 32'h00000493;
          45:    rdata = 32'h00000513;
          46:    rdata = 32'h00000593;
          47:    rdata = 32'h00000613;
          48:    rdata = 32'h00000693;
          49:    rdata = 32'h00000713;
          50:    rdata = 32'h00000793;
          51:    rdata = 32'h00000813;
          52:    rdata = 32'h00000893;
          53:    rdata = 32'h00000913;
          54:    rdata = 32'h00000993;
          55:    rdata = 32'h00000a13;
          56:    rdata = 32'h00000a93;
          57:    rdata = 32'h00000b13;
          58:    rdata = 32'h00000b93;
          59:    rdata = 32'h00000c13;
          60:    rdata = 32'h00000c93;
          61:    rdata = 32'h00000d13;
          62:    rdata = 32'h00000d93;
          63:    rdata = 32'h00000e13;
          64:    rdata = 32'h00000e93;
          65:    rdata = 32'h00000f13;
          66:    rdata = 32'h00000f93;
          67:    rdata = 32'h000f4117;
          68:    rdata = 32'hef410113;
          69:    rdata = 32'h000f0297;
          70:    rdata = 32'heec28293;
          71:    rdata = 32'h000f0317;
          72:    rdata = 32'hf5830313;
          73:    rdata = 32'h0062d863;
          74:    rdata = 32'h0002a023;
          75:    rdata = 32'h00428293;
          76:    rdata = 32'hfe535ce3;
          77:    rdata = 32'h00001297;
          78:    rdata = 32'h3f428293;
          79:    rdata = 32'h000f0317;
          80:    rdata = 32'hec430313;
          81:    rdata = 32'h000f0397;
          82:    rdata = 32'hebc38393;
          83:    rdata = 32'h00735c63;
          84:    rdata = 32'h0002ae03;
          85:    rdata = 32'h01c32023;
          86:    rdata = 32'h00428293;
          87:    rdata = 32'h00430313;
          88:    rdata = 32'hfe7348e3;
          89:    rdata = 32'h00001297;
          90:    rdata = 32'h1b828293;
          91:    rdata = 32'h00001317;
          92:    rdata = 32'h1c030313;
          93:    rdata = 32'h0062da63;
          94:    rdata = 32'h0002a783;
          95:    rdata = 32'h000780e7;
          96:    rdata = 32'h00428293;
          97:    rdata = 32'hfe62cae3;
          98:    rdata = 32'h00000513;
          99:    rdata = 32'h00000593;
         100:    rdata = 32'h118010ef;
         101:    rdata = 32'hdca27119;
         102:    rdata = 32'h00001597;
         103:    rdata = 32'h24058593;
         104:    rdata = 32'h0517842a;
         105:    rdata = 32'h0513000f;
         106:    rdata = 32'hde86eaa5;
         107:    rdata = 32'h549000ef;
         108:    rdata = 32'h0613006c;
         109:    rdata = 32'h05170640;
         110:    rdata = 32'h0513000f;
         111:    rdata = 32'h00efe965;
         112:    rdata = 32'h006c4d70;
         113:    rdata = 32'h227d8522;
         114:    rdata = 32'h546650f6;
         115:    rdata = 32'h80826109;
         116:    rdata = 32'h00001597;
         117:    rdata = 32'h20c58593;
         118:    rdata = 32'h000f0517;
         119:    rdata = 32'he7450513;
         120:    rdata = 32'h5150006f;
         121:    rdata = 32'h15171141;
         122:    rdata = 32'h05130000;
         123:    rdata = 32'hc6062865;
         124:    rdata = 32'h00efc422;
         125:    rdata = 32'h842a10b0;
         126:    rdata = 32'h00001517;
         127:    rdata = 32'h27850513;
         128:    rdata = 32'h0fd000ef;
         129:    rdata = 32'h0ff47593;
         130:    rdata = 32'h40b24422;
         131:    rdata = 32'h00a03633;
         132:    rdata = 32'h000f0517;
         133:    rdata = 32'hdf050513;
         134:    rdata = 32'h006f0141;
         135:    rdata = 32'h11012690;
         136:    rdata = 32'hcc22ce06;
         137:    rdata = 32'h0113ca26;
         138:    rdata = 32'h06138101;
         139:    rdata = 32'h45810400;
         140:    rdata = 32'h00ef850a;
         141:    rdata = 32'h858a61f0;
         142:    rdata = 32'h000f0517;
         143:    rdata = 32'hde850513;
         144:    rdata = 32'h2bb000ef;
         145:    rdata = 32'h000f0517;
         146:    rdata = 32'he2050513;
         147:    rdata = 32'h10d000ef;
         148:    rdata = 32'h0597842a;
         149:    rdata = 32'h8593000f;
         150:    rdata = 32'h850ae0e5;
         151:    rdata = 32'h05172695;
         152:    rdata = 32'h0513000f;
         153:    rdata = 32'h00efe065;
         154:    rdata = 32'h05b30f30;
         155:    rdata = 32'h15174085;
         156:    rdata = 32'h05130000;
         157:    rdata = 32'h22fd20a5;
         158:    rdata = 32'h0084840a;
         159:    rdata = 32'h7c045503;
         160:    rdata = 32'h22710409;
         161:    rdata = 32'hfe941ce3;
         162:    rdata = 32'h7f010113;
         163:    rdata = 32'h446240f2;
         164:    rdata = 32'h610544d2;
         165:    rdata = 32'h715d8082;
         166:    rdata = 32'h04000593;
         167:    rdata = 32'h000f0517;
         168:    rdata = 32'hd8450513;
         169:    rdata = 32'hc4a2c686;
         170:    rdata = 32'h281000ef;
         171:    rdata = 32'h04000613;
         172:    rdata = 32'h850a4581;
         173:    rdata = 32'h59d000ef;
         174:    rdata = 32'h0517858a;
         175:    rdata = 32'h0513000f;
         176:    rdata = 32'h00efd665;
         177:    rdata = 32'h05172390;
         178:    rdata = 32'h0513000f;
         179:    rdata = 32'h00efd9e5;
         180:    rdata = 32'h842a08b0;
         181:    rdata = 32'h000f0517;
         182:    rdata = 32'hd8c50513;
         183:    rdata = 32'h0517292d;
         184:    rdata = 32'h0513000f;
         185:    rdata = 32'h00efd865;
         186:    rdata = 32'h04330730;
         187:    rdata = 32'h15974085;
         188:    rdata = 32'h85930000;
         189:    rdata = 32'h051719a5;
         190:    rdata = 32'h0513000f;
         191:    rdata = 32'h00efd565;
         192:    rdata = 32'h85a23f70;
         193:    rdata = 32'h40b64426;
         194:    rdata = 32'h00001517;
         195:    rdata = 32'h19c50513;
         196:    rdata = 32'haa896161;
         197:    rdata = 32'hcc221101;
         198:    rdata = 32'hc84aca26;
         199:    rdata = 32'hc452c64e;
         200:    rdata = 32'h842ace06;
         201:    rdata = 32'h14974a11;
         202:    rdata = 32'h84930000;
         203:    rdata = 32'h19970064;
         204:    rdata = 32'h89930000;
         205:    rdata = 32'h091718a9;
         206:    rdata = 32'h0913000f;
         207:    rdata = 32'h8522d169;
         208:    rdata = 32'h6ee33d91;
         209:    rdata = 32'h1793feaa;
         210:    rdata = 32'h97a60025;
         211:    rdata = 32'h97a6439c;
         212:    rdata = 32'h85228782;
         213:    rdata = 32'hb7e53db5;
         214:    rdata = 32'h35698522;
         215:    rdata = 32'h8522b7cd;
         216:    rdata = 32'hbff13d7d;
         217:    rdata = 32'h3f058522;
         218:    rdata = 32'h85cebfd9;
         219:    rdata = 32'h00ef854a;
         220:    rdata = 32'hb7f13870;
         221:    rdata = 32'hc4221141;
         222:    rdata = 32'h8522842e;
         223:    rdata = 32'h00001597;
         224:    rdata = 32'h15458593;
         225:    rdata = 32'h00efc606;
         226:    rdata = 32'h87aa5a70;
         227:    rdata = 32'h1597cd0d;
         228:    rdata = 32'h85930000;
         229:    rdata = 32'h852214a5;
         230:    rdata = 32'h595000ef;
         231:    rdata = 32'hc5054785;
         232:    rdata = 32'h00001597;
         233:    rdata = 32'h14058593;
         234:    rdata = 32'h00ef8522;
         235:    rdata = 32'h47895830;
         236:    rdata = 32'h1597c919;
         237:    rdata = 32'h85930000;
         238:    rdata = 32'h852213a5;
         239:    rdata = 32'h571000ef;
         240:    rdata = 32'h00a037b3;
         241:    rdata = 32'h40b2078d;
         242:    rdata = 32'h853e4422;
         243:    rdata = 32'h80820141;
         244:    rdata = 32'h85aa7119;
         245:    rdata = 32'hde860068;
         246:    rdata = 32'h15972b61;
         247:    rdata = 32'h85930000;
         248:    rdata = 32'h00680f25;
         249:    rdata = 32'h006c2b79;
         250:    rdata = 32'h000f0517;
         251:    rdata = 32'hc6450513;
         252:    rdata = 32'h305000ef;
         253:    rdata = 32'h610950f6;
         254:    rdata = 32'h11018082;
         255:    rdata = 32'h004885aa;
         256:    rdata = 32'h2525ce06;
         257:    rdata = 32'h37e90048;
         258:    rdata = 32'h610540f2;
         259:    rdata = 32'h11018082;
         260:    rdata = 32'h004885aa;
         261:    rdata = 32'h2569ce06;
         262:    rdata = 32'h3f5d0048;
         263:    rdata = 32'h610540f2;
         264:    rdata = 32'h71198082;
         265:    rdata = 32'h842edca2;
         266:    rdata = 32'h006885aa;
         267:    rdata = 32'h2389de86;
         268:    rdata = 32'h00001597;
         269:    rdata = 32'h0d058593;
         270:    rdata = 32'h23a10068;
         271:    rdata = 32'h006885a2;
         272:    rdata = 32'h15972389;
         273:    rdata = 32'h85930000;
         274:    rdata = 32'h006808a5;
         275:    rdata = 32'h006c2b1d;
         276:    rdata = 32'h000f0517;
         277:    rdata = 32'hbfc50513;
         278:    rdata = 32'h29d000ef;
         279:    rdata = 32'h546650f6;
         280:    rdata = 32'h80826109;
         281:    rdata = 32'hcc221101;
         282:    rdata = 32'h0048842a;
         283:    rdata = 32'h2b75ce06;
         284:    rdata = 32'h8522004c;
         285:    rdata = 32'h40f2377d;
         286:    rdata = 32'h61054462;
         287:    rdata = 32'h11018082;
         288:    rdata = 32'h842acc22;
         289:    rdata = 32'hce060048;
         290:    rdata = 32'h004c2d21;
         291:    rdata = 32'h3f518522;
         292:    rdata = 32'h446240f2;
         293:    rdata = 32'h80826105;
         294:    rdata = 32'hdaa67119;
         295:    rdata = 32'h85aa84ae;
         296:    rdata = 32'hde860068;
         297:    rdata = 32'h8432dca2;
         298:    rdata = 32'h159721e1;
         299:    rdata = 32'h85930000;
         300:    rdata = 32'h006805a5;
         301:    rdata = 32'h85a621f9;
         302:    rdata = 32'h21e10068;
         303:    rdata = 32'h00001597;
         304:    rdata = 32'h04c58593;
         305:    rdata = 32'h29750068;
         306:    rdata = 32'h006885a2;
         307:    rdata = 32'h1597295d;
         308:    rdata = 32'h85930000;
         309:    rdata = 32'h0068ffe5;
         310:    rdata = 32'h006c216d;
         311:    rdata = 32'h000f0517;
         312:    rdata = 32'hb7050513;
         313:    rdata = 32'h211000ef;
         314:    rdata = 32'h546650f6;
         315:    rdata = 32'h610954d6;
         316:    rdata = 32'h71798082;
         317:    rdata = 32'h842ad422;
         318:    rdata = 32'hd6060028;
         319:    rdata = 32'h84b2d226;
         320:    rdata = 32'h85a62345;
         321:    rdata = 32'h23150848;
         322:    rdata = 32'h002c0850;
         323:    rdata = 32'h37698522;
         324:    rdata = 32'h542250b2;
         325:    rdata = 32'h61455492;
         326:    rdata = 32'h71798082;
         327:    rdata = 32'h842ad422;
         328:    rdata = 32'hd6060028;
         329:    rdata = 32'h84b2d226;
         330:    rdata = 32'h85a62ba5;
         331:    rdata = 32'h2b8d0848;
         332:    rdata = 32'h002c0850;
         333:    rdata = 32'h378d8522;
         334:    rdata = 32'h542250b2;
         335:    rdata = 32'h61455492;
         336:    rdata = 32'h11018082;
         337:    rdata = 32'h842acc22;
         338:    rdata = 32'h000f0517;
         339:    rdata = 32'haf450513;
         340:    rdata = 32'hca26ce06;
         341:    rdata = 32'hc64ec84a;
         342:    rdata = 32'h00efc452;
         343:    rdata = 32'h05170d70;
         344:    rdata = 32'h0513000f;
         345:    rdata = 32'h00efade5;
         346:    rdata = 32'h04977ec0;
         347:    rdata = 32'h8493000f;
         348:    rdata = 32'h8526ad24;
         349:    rdata = 32'h7ea000ef;
         350:    rdata = 32'h44fddd6d;
         351:    rdata = 32'h000f0917;
         352:    rdata = 32'hac090913;
         353:    rdata = 32'h000f0a17;
         354:    rdata = 32'ha9ca0a13;
         355:    rdata = 32'h854a59fd;
         356:    rdata = 32'h7c2000ef;
         357:    rdata = 32'h00ef854a;
         358:    rdata = 32'hdd6d7c80;
         359:    rdata = 32'h00649593;
         360:    rdata = 32'h855295a2;
         361:    rdata = 32'h00ef14fd;
         362:    rdata = 32'h92e375c0;
         363:    rdata = 32'h40f2ff34;
         364:    rdata = 32'h44628522;
         365:    rdata = 32'h494244d2;
         366:    rdata = 32'h4a2249b2;
         367:    rdata = 32'h80826105;
         368:    rdata = 32'hcc221101;
         369:    rdata = 32'h0517842a;
         370:    rdata = 32'h0513000f;
         371:    rdata = 32'hce06a765;
         372:    rdata = 32'h00efc62e;
         373:    rdata = 32'h05170790;
         374:    rdata = 32'h0513000f;
         375:    rdata = 32'h00efa665;
         376:    rdata = 32'h45b27740;
         377:    rdata = 32'h3fb18522;
         378:    rdata = 32'h852240f2;
         379:    rdata = 32'h61054462;
         380:    rdata = 32'h715d8082;
         381:    rdata = 32'h872e878a;
         382:    rdata = 32'hc4a2c686;
         383:    rdata = 32'h85bec2a6;
         384:    rdata = 32'h00e79023;
         385:    rdata = 32'h07890094;
         386:    rdata = 32'hfed79ce3;
         387:    rdata = 32'h000f0517;
         388:    rdata = 32'ha1450513;
         389:    rdata = 32'h051725dd;
         390:    rdata = 32'h0513000f;
         391:    rdata = 32'h00efa265;
         392:    rdata = 32'h05170130;
         393:    rdata = 32'h0513000f;
         394:    rdata = 32'h00efa1a5;
         395:    rdata = 32'h04177280;
         396:    rdata = 32'h0413000f;
         397:    rdata = 32'h8522a0e4;
         398:    rdata = 32'h726000ef;
         399:    rdata = 32'h0413dd6d;
         400:    rdata = 32'h04970200;
         401:    rdata = 32'h8493000f;
         402:    rdata = 32'h85269fa4;
         403:    rdata = 32'h706000ef;
         404:    rdata = 32'h00ef8526;
         405:    rdata = 32'hdd6d70c0;
         406:    rdata = 32'hf865147d;
         407:    rdata = 32'h442640b6;
         408:    rdata = 32'h61614496;
         409:    rdata = 32'h11418082;
         410:    rdata = 32'h3761c606;
         411:    rdata = 32'h000f0517;
         412:    rdata = 32'h9d050513;
         413:    rdata = 32'h7ca000ef;
         414:    rdata = 32'h051740b2;
         415:    rdata = 32'h0513000f;
         416:    rdata = 32'h01419c25;
         417:    rdata = 32'h1101a5f9;
         418:    rdata = 32'h000f0517;
         419:    rdata = 32'h9b450513;
         420:    rdata = 32'hcc22ce06;
         421:    rdata = 32'hc84aca26;
         422:    rdata = 32'hc64e84ae;
         423:    rdata = 32'h794000ef;
         424:    rdata = 32'h000f0517;
         425:    rdata = 32'h99c50513;
         426:    rdata = 32'h0417256d;
         427:    rdata = 32'h0413000f;
         428:    rdata = 32'h85229924;
         429:    rdata = 32'hdd75256d;
         430:    rdata = 32'h7c048413;
         431:    rdata = 32'h000f0997;
         432:    rdata = 32'h96498993;
         433:    rdata = 32'h000f0917;
         434:    rdata = 32'h97890913;
         435:    rdata = 32'h85a2854e;
         436:    rdata = 32'h854a252d;
         437:    rdata = 32'h854a2dbd;
         438:    rdata = 32'hdd752559;
         439:    rdata = 32'hfc040793;
         440:    rdata = 32'h00849963;
         441:    rdata = 32'h446240f2;
         442:    rdata = 32'h494244d2;
         443:    rdata = 32'h610549b2;
         444:    rdata = 32'h843e8082;
         445:    rdata = 32'h1141bfe1;
         446:    rdata = 32'h3771c606;
         447:    rdata = 32'h000f0517;
         448:    rdata = 32'h94050513;
         449:    rdata = 32'h73a000ef;
         450:    rdata = 32'h051740b2;
         451:    rdata = 32'h0513000f;
         452:    rdata = 32'h01419325;
         453:    rdata = 32'h7139ad3d;
         454:    rdata = 32'hd452737d;
         455:    rdata = 32'h81030313;
         456:    rdata = 32'hdc226a09;
         457:    rdata = 32'hd84ada26;
         458:    rdata = 32'hd256d64e;
         459:    rdata = 32'hce5ed05a;
         460:    rdata = 32'hde06cc62;
         461:    rdata = 32'h800a0793;
         462:    rdata = 32'h978a911a;
         463:    rdata = 32'h84b3747d;
         464:    rdata = 32'h892a0087;
         465:    rdata = 32'h45816605;
         466:    rdata = 32'h00ef8526;
         467:    rdata = 32'h07931070;
         468:    rdata = 32'h0413800a;
         469:    rdata = 32'h978a8004;
         470:    rdata = 32'h943e6a05;
         471:    rdata = 32'h880a0a13;
         472:    rdata = 32'h89934b01;
         473:    rdata = 32'h0b938004;
         474:    rdata = 32'h8aa60804;
         475:    rdata = 32'h0c139a22;
         476:    rdata = 32'h854a0800;
         477:    rdata = 32'h080b4433;
         478:    rdata = 32'h35f585a2;
         479:    rdata = 32'h85ca854e;
         480:    rdata = 32'h855e3581;
         481:    rdata = 32'h0e138826;
         482:    rdata = 32'h0693f805;
         483:    rdata = 32'h03131808;
         484:    rdata = 32'h07130405;
         485:    rdata = 32'h07931008;
         486:    rdata = 32'h05930808;
         487:    rdata = 32'h88aafc05;
         488:    rdata = 32'h5e838642;
         489:    rdata = 32'h5f03000e;
         490:    rdata = 32'h76630026;
         491:    rdata = 32'h102301df;
         492:    rdata = 32'h11230086;
         493:    rdata = 32'h5e8301d6;
         494:    rdata = 32'h5f03002e;
         495:    rdata = 32'h76630066;
         496:    rdata = 32'h122301df;
         497:    rdata = 32'h13230086;
         498:    rdata = 32'h5e8301d6;
         499:    rdata = 32'h5f03004e;
         500:    rdata = 32'h766300a6;
         501:    rdata = 32'h142301df;
         502:    rdata = 32'h15230086;
         503:    rdata = 32'h5e8301d6;
         504:    rdata = 32'h5f03006e;
         505:    rdata = 32'h766300e6;
         506:    rdata = 32'h162301df;
         507:    rdata = 32'h17230086;
         508:    rdata = 32'hde8301d6;
         509:    rdata = 32'hdf030005;
         510:    rdata = 32'h76630027;
         511:    rdata = 32'h902301df;
         512:    rdata = 32'h91230087;
         513:    rdata = 32'hde8301d7;
         514:    rdata = 32'hdf030025;
         515:    rdata = 32'h76630067;
         516:    rdata = 32'h922301df;
         517:    rdata = 32'h93230087;
         518:    rdata = 32'hde8301d7;
         519:    rdata = 32'hdf030045;
         520:    rdata = 32'h766300a7;
         521:    rdata = 32'h942301df;
         522:    rdata = 32'h95230087;
         523:    rdata = 32'hde8301d7;
         524:    rdata = 32'hdf030065;
         525:    rdata = 32'h766300e7;
         526:    rdata = 32'h962301df;
         527:    rdata = 32'h97230087;
         528:    rdata = 32'hde8301d7;
         529:    rdata = 32'h5f030008;
         530:    rdata = 32'h76630027;
         531:    rdata = 32'h102301df;
         532:    rdata = 32'h11230087;
         533:    rdata = 32'hde8301d7;
         534:    rdata = 32'h5f030028;
         535:    rdata = 32'h76630067;
         536:    rdata = 32'h122301df;
         537:    rdata = 32'h13230087;
         538:    rdata = 32'hde8301d7;
         539:    rdata = 32'h5f030048;
         540:    rdata = 32'h766300a7;
         541:    rdata = 32'h142301df;
         542:    rdata = 32'h15230087;
         543:    rdata = 32'hde8301d7;
         544:    rdata = 32'h5f030068;
         545:    rdata = 32'h766300e7;
         546:    rdata = 32'h162301df;
         547:    rdata = 32'h17230087;
         548:    rdata = 32'h5e8301d7;
         549:    rdata = 32'hdf030003;
         550:    rdata = 32'h76630026;
         551:    rdata = 32'h902301df;
         552:    rdata = 32'h91230086;
         553:    rdata = 32'h5e8301d6;
         554:    rdata = 32'hdf030023;
         555:    rdata = 32'h76630066;
         556:    rdata = 32'h922301df;
         557:    rdata = 32'h93230086;
         558:    rdata = 32'h5e8301d6;
         559:    rdata = 32'hdf030043;
         560:    rdata = 32'h766300a6;
         561:    rdata = 32'h942301df;
         562:    rdata = 32'h95230086;
         563:    rdata = 32'h5e8301d6;
         564:    rdata = 32'hdf030063;
         565:    rdata = 32'h766300e6;
         566:    rdata = 32'h962301df;
         567:    rdata = 32'h97230086;
         568:    rdata = 32'h05a101d6;
         569:    rdata = 32'h06410e21;
         570:    rdata = 32'h032106c1;
         571:    rdata = 32'h08a10741;
         572:    rdata = 32'h98e307c1;
         573:    rdata = 32'h8513eaa5;
         574:    rdata = 32'h08131005;
         575:    rdata = 32'h14e32008;
         576:    rdata = 32'h0b05e945;
         577:    rdata = 32'he78b17e3;
         578:    rdata = 32'h777d6789;
         579:    rdata = 32'h80078793;
         580:    rdata = 32'h0713978a;
         581:    rdata = 32'h973e8007;
         582:    rdata = 32'h94be6785;
         583:    rdata = 32'h86ba87d6;
         584:    rdata = 32'h080a8a93;
         585:    rdata = 32'h0007d603;
         586:    rdata = 32'h06890791;
         587:    rdata = 32'hfec69f23;
         588:    rdata = 32'hfefa9ae3;
         589:    rdata = 32'h04070713;
         590:    rdata = 32'hfe9a92e3;
         591:    rdata = 32'h75fd6789;
         592:    rdata = 32'h80078793;
         593:    rdata = 32'h8593978a;
         594:    rdata = 32'h854a8005;
         595:    rdata = 32'h336595be;
         596:    rdata = 32'h03136305;
         597:    rdata = 32'h911a7f03;
         598:    rdata = 32'h546250f2;
         599:    rdata = 32'h594254d2;
         600:    rdata = 32'h5a2259b2;
         601:    rdata = 32'h5b025a92;
         602:    rdata = 32'h4c624bf2;
         603:    rdata = 32'h80826121;
         604:    rdata = 32'hc70387aa;
         605:    rdata = 32'h05850005;
         606:    rdata = 32'h8fa30785;
         607:    rdata = 32'hfb75fee7;
         608:    rdata = 32'h87aa8082;
         609:    rdata = 32'h0007c683;
         610:    rdata = 32'h0785873e;
         611:    rdata = 32'hc783fee5;
         612:    rdata = 32'h05850005;
         613:    rdata = 32'h0fa30705;
         614:    rdata = 32'hfbf5fef7;
         615:    rdata = 32'h47838082;
         616:    rdata = 32'hc7030005;
         617:    rdata = 32'h87630005;
         618:    rdata = 32'h557d00e7;
         619:    rdata = 32'h00e7e963;
         620:    rdata = 32'h80824505;
         621:    rdata = 32'h0505c781;
         622:    rdata = 32'hb7d50585;
         623:    rdata = 32'h80824501;
         624:    rdata = 32'h450187aa;
         625:    rdata = 32'h00a78733;
         626:    rdata = 32'h00074703;
         627:    rdata = 32'h0505c319;
         628:    rdata = 32'h8082bfd5;
         629:    rdata = 32'h0c634789;
         630:    rdata = 32'h479102f6;
         631:    rdata = 32'h02f60d63;
         632:    rdata = 32'h47814705;
         633:    rdata = 32'h00e61463;
         634:    rdata = 32'h06400793;
         635:    rdata = 32'hcb8d4629;
         636:    rdata = 32'h02f5d733;
         637:    rdata = 32'h76930505;
         638:    rdata = 32'h86b30ff7;
         639:    rdata = 32'h071302f6;
         640:    rdata = 32'h0fa30307;
         641:    rdata = 32'hd7b3fee5;
         642:    rdata = 32'h8d9502c7;
         643:    rdata = 32'h6789b7cd;
         644:    rdata = 32'h71078793;
         645:    rdata = 32'hd7b7bfe1;
         646:    rdata = 32'h87933b9a;
         647:    rdata = 32'hb7f9a007;
         648:    rdata = 32'h00050023;
         649:    rdata = 32'h46058082;
         650:    rdata = 32'h1101b775;
         651:    rdata = 32'h4611cc22;
         652:    rdata = 32'h0048842a;
         653:    rdata = 32'h3f79ce06;
         654:    rdata = 32'h0713004c;
         655:    rdata = 32'hc7830300;
         656:    rdata = 32'h94630005;
         657:    rdata = 32'h058500e7;
         658:    rdata = 32'he391bfdd;
         659:    rdata = 32'h852215fd;
         660:    rdata = 32'h40f23705;
         661:    rdata = 32'h61054462;
         662:    rdata = 32'h07938082;
         663:    rdata = 32'h06060300;
         664:    rdata = 32'h0ff67613;
         665:    rdata = 32'h00f50023;
         666:    rdata = 32'h07800793;
         667:    rdata = 32'h00f500a3;
         668:    rdata = 32'h87b24825;
         669:    rdata = 32'hf713c385;
         670:    rdata = 32'h069300f5;
         671:    rdata = 32'h64630577;
         672:    rdata = 32'h069300e8;
         673:    rdata = 32'h07330307;
         674:    rdata = 32'h00a300f5;
         675:    rdata = 32'h819100d7;
         676:    rdata = 32'hb7cd17fd;
         677:    rdata = 32'h01239532;
         678:    rdata = 32'h80820005;
         679:    rdata = 32'hbf754605;
         680:    rdata = 32'hbf654611;
         681:    rdata = 32'h47834725;
         682:    rdata = 32'h87930005;
         683:    rdata = 32'hf793fd07;
         684:    rdata = 32'h68630ff7;
         685:    rdata = 32'h478300f7;
         686:    rdata = 32'h05050015;
         687:    rdata = 32'h4505f7ed;
         688:    rdata = 32'h45018082;
         689:    rdata = 32'h46038082;
         690:    rdata = 32'h07130005;
         691:    rdata = 32'h87aa02d0;
         692:    rdata = 32'h15634681;
         693:    rdata = 32'h079300e6;
         694:    rdata = 32'h46850015;
         695:    rdata = 32'h46294501;
         696:    rdata = 32'h0007c703;
         697:    rdata = 32'h0533cb01;
         698:    rdata = 32'h071302c5;
         699:    rdata = 32'h0785fd07;
         700:    rdata = 32'hb7fd953a;
         701:    rdata = 32'h0533c299;
         702:    rdata = 32'h808240a0;
         703:    rdata = 32'hc5227175;
         704:    rdata = 32'hc14ac326;
         705:    rdata = 32'hc706dece;
         706:    rdata = 32'hf41784aa;
         707:    rdata = 32'h0413000e;
         708:    rdata = 32'h19975424;
         709:    rdata = 32'h89930000;
         710:    rdata = 32'h19179ee9;
         711:    rdata = 32'h09130000;
         712:    rdata = 32'h85a69f29;
         713:    rdata = 32'h26f98522;
         714:    rdata = 32'h852285ce;
         715:    rdata = 32'h061326e1;
         716:    rdata = 32'h006c0640;
         717:    rdata = 32'h2eb98522;
         718:    rdata = 32'h37ad0068;
         719:    rdata = 32'h85cae509;
         720:    rdata = 32'h2e4d8522;
         721:    rdata = 32'h0068bff9;
         722:    rdata = 32'h40ba3fbd;
         723:    rdata = 32'h449a442a;
         724:    rdata = 32'h59f6490a;
         725:    rdata = 32'h80826149;
         726:    rdata = 32'hb0002573;
         727:    rdata = 32'hb80025f3;
         728:    rdata = 32'h00018082;
         729:    rdata = 32'h00010001;
         730:    rdata = 32'h00010001;
         731:    rdata = 32'h15fd0001;
         732:    rdata = 32'h8082f9ed;
         733:    rdata = 32'h300462f3;
         734:    rdata = 32'hc10c8082;
         735:    rdata = 32'ha2f362c1;
         736:    rdata = 32'h80823042;
         737:    rdata = 32'h02b7c14c;
         738:    rdata = 32'ha2f30002;
         739:    rdata = 32'h80823042;
         740:    rdata = 32'hcc3e7139;
         741:    rdata = 32'hdc16de06;
         742:    rdata = 32'hd81eda1a;
         743:    rdata = 32'hd42ed62a;
         744:    rdata = 32'hd036d232;
         745:    rdata = 32'hca42ce3a;
         746:    rdata = 32'hc672c846;
         747:    rdata = 32'hc27ac476;
         748:    rdata = 32'hf797c07e;
         749:    rdata = 32'ha783000e;
         750:    rdata = 32'h97824b27;
         751:    rdata = 32'h52e250f2;
         752:    rdata = 32'h53c25352;
         753:    rdata = 32'h55a25532;
         754:    rdata = 32'h56825612;
         755:    rdata = 32'h47e24772;
         756:    rdata = 32'h48c24852;
         757:    rdata = 32'h4ea24e32;
         758:    rdata = 32'h4f824f12;
         759:    rdata = 32'h00736121;
         760:    rdata = 32'h71393020;
         761:    rdata = 32'hde06cc3e;
         762:    rdata = 32'hda1adc16;
         763:    rdata = 32'hd62ad81e;
         764:    rdata = 32'hd232d42e;
         765:    rdata = 32'hce3ad036;
         766:    rdata = 32'hc846ca42;
         767:    rdata = 32'hc476c672;
         768:    rdata = 32'hc07ec27a;
         769:    rdata = 32'h000ef797;
         770:    rdata = 32'h4647a783;
         771:    rdata = 32'h50f29782;
         772:    rdata = 32'h535252e2;
         773:    rdata = 32'h553253c2;
         774:    rdata = 32'h561255a2;
         775:    rdata = 32'h47725682;
         776:    rdata = 32'h485247e2;
         777:    rdata = 32'h4e3248c2;
         778:    rdata = 32'h4f124ea2;
         779:    rdata = 32'h61214f82;
         780:    rdata = 32'h30200073;
         781:    rdata = 32'h00458793;
         782:    rdata = 32'h8793c15c;
         783:    rdata = 32'hc51c0085;
         784:    rdata = 32'h00c58793;
         785:    rdata = 32'h8793c55c;
         786:    rdata = 32'hc91c0105;
         787:    rdata = 32'h01458793;
         788:    rdata = 32'hc95cc10c;
         789:    rdata = 32'h01858793;
         790:    rdata = 32'hcd1c05f1;
         791:    rdata = 32'h8082cd4c;
         792:    rdata = 32'h4388455c;
         793:    rdata = 32'h97b34785;
         794:    rdata = 32'h8d7d00b7;
         795:    rdata = 32'h00a03533;
         796:    rdata = 32'h451c8082;
         797:    rdata = 32'h8e3d439c;
         798:    rdata = 32'h8e3d8e6d;
         799:    rdata = 32'hc390451c;
         800:    rdata = 32'h47858082;
         801:    rdata = 32'h00b61633;
         802:    rdata = 32'h00b795b3;
         803:    rdata = 32'h1141b7dd;
         804:    rdata = 32'hc226c422;
         805:    rdata = 32'h842ac606;
         806:    rdata = 32'h37d984ae;
         807:    rdata = 32'h00154613;
         808:    rdata = 32'h44228522;
         809:    rdata = 32'h85a640b2;
         810:    rdata = 32'h76134492;
         811:    rdata = 32'h01410ff6;
         812:    rdata = 32'h455cbfc9;
         813:    rdata = 32'h55134388;
         814:    rdata = 32'h80824915;
         815:    rdata = 32'h4388455c;
         816:    rdata = 32'h49055513;
         817:    rdata = 32'h862e8082;
         818:    rdata = 32'hbf6545bd;
         819:    rdata = 32'h00858713;
         820:    rdata = 32'h05058793;
         821:    rdata = 32'hc91cc518;
         822:    rdata = 32'h01058713;
         823:    rdata = 32'h010107b7;
         824:    rdata = 32'h8613c558;
         825:    rdata = 32'h87130045;
         826:    rdata = 32'h87931007;
         827:    rdata = 32'hc10c2007;
         828:    rdata = 32'hc958c150;
         829:    rdata = 32'h0571cd1c;
         830:    rdata = 32'h4548a81d;
         831:    rdata = 32'h04000613;
         832:    rdata = 32'h87aaac15;
         833:    rdata = 32'h4b8c852e;
         834:    rdata = 32'h04000613;
         835:    rdata = 32'h495ca425;
         836:    rdata = 32'hc3984198;
         837:    rdata = 32'h41d8495c;
         838:    rdata = 32'h4598c3d8;
         839:    rdata = 32'hc798495c;
         840:    rdata = 32'h495c45d8;
         841:    rdata = 32'h8082c7d8;
         842:    rdata = 32'hc38c4d1c;
         843:    rdata = 32'hc10c8082;
         844:    rdata = 32'h15b7c150;
         845:    rdata = 32'h06130101;
         846:    rdata = 32'h05214000;
         847:    rdata = 32'h4118a2dd;
         848:    rdata = 32'h0015c593;
         849:    rdata = 32'h0015f793;
         850:    rdata = 32'h99f9430c;
         851:    rdata = 32'hc30c8ddd;
         852:    rdata = 32'h41188082;
         853:    rdata = 32'he793431c;
         854:    rdata = 32'hc31c0027;
         855:    rdata = 32'h415c8082;
         856:    rdata = 32'h89054388;
         857:    rdata = 32'h71398082;
         858:    rdata = 32'h4411dc22;
         859:    rdata = 32'h02864433;
         860:    rdata = 32'hda264118;
         861:    rdata = 32'hd64ed84a;
         862:    rdata = 32'hd256d452;
         863:    rdata = 32'hcc62ce5e;
         864:    rdata = 32'hd05ade06;
         865:    rdata = 32'h84aa431c;
         866:    rdata = 32'h9bf989ae;
         867:    rdata = 32'hc31c8932;
         868:    rdata = 32'h4a814a01;
         869:    rdata = 32'h0b934c11;
         870:    rdata = 32'hd9630085;
         871:    rdata = 32'h4781028a;
         872:    rdata = 32'h01498633;
         873:    rdata = 32'h00f606b3;
         874:    rdata = 32'h0006c683;
         875:    rdata = 32'h973e0078;
         876:    rdata = 32'h00d70023;
         877:    rdata = 32'h97e30785;
         878:    rdata = 32'h4b32ff87;
         879:    rdata = 32'h855e85d2;
         880:    rdata = 32'h202322a5;
         881:    rdata = 32'h0a850165;
         882:    rdata = 32'hbfc10a11;
         883:    rdata = 32'h54334581;
         884:    rdata = 32'h15930ab4;
         885:    rdata = 32'h05330024;
         886:    rdata = 32'h0a6340b9;
         887:    rdata = 32'h478102b9;
         888:    rdata = 32'h4701468d;
         889:    rdata = 32'h00a7d763;
         890:    rdata = 32'h00f58733;
         891:    rdata = 32'h4703974e;
         892:    rdata = 32'h00700007;
         893:    rdata = 32'h0023963e;
         894:    rdata = 32'h078500e6;
         895:    rdata = 32'hfed793e3;
         896:    rdata = 32'h000107a3;
         897:    rdata = 32'h85134432;
         898:    rdata = 32'h2a390084;
         899:    rdata = 32'h4098c100;
         900:    rdata = 32'he793431c;
         901:    rdata = 32'hc31c0017;
         902:    rdata = 32'h546250f2;
         903:    rdata = 32'h594254d2;
         904:    rdata = 32'h5a2259b2;
         905:    rdata = 32'h5b025a92;
         906:    rdata = 32'h4c624bf2;
         907:    rdata = 32'h80826121;
         908:    rdata = 32'h06700613;
         909:    rdata = 32'h00000597;
         910:    rdata = 32'h50c58593;
         911:    rdata = 32'h4625b72d;
         912:    rdata = 32'h00000597;
         913:    rdata = 32'h56858593;
         914:    rdata = 32'h4625bf39;
         915:    rdata = 32'h00000597;
         916:    rdata = 32'h56858593;
         917:    rdata = 32'h8793bf09;
         918:    rdata = 32'hc15c0045;
         919:    rdata = 32'h00858793;
         920:    rdata = 32'h8793c51c;
         921:    rdata = 32'hc55c00c5;
         922:    rdata = 32'h01058793;
         923:    rdata = 32'h4799c91c;
         924:    rdata = 32'h8823c10c;
         925:    rdata = 32'h419c00f5;
         926:    rdata = 32'h0017e793;
         927:    rdata = 32'h8082c19c;
         928:    rdata = 32'h439c415c;
         929:    rdata = 32'hdfed8b85;
         930:    rdata = 32'hc503455c;
         931:    rdata = 32'h75130007;
         932:    rdata = 32'h80820ff5;
         933:    rdata = 32'hcc221101;
         934:    rdata = 32'hc84aca26;
         935:    rdata = 32'hc256c64e;
         936:    rdata = 32'hc452ce06;
         937:    rdata = 32'h892e84aa;
         938:    rdata = 32'h440189b2;
         939:    rdata = 32'h58634aa9;
         940:    rdata = 32'h85260334;
         941:    rdata = 32'h00890a33;
         942:    rdata = 32'h002337e1;
         943:    rdata = 32'h1e6300aa;
         944:    rdata = 32'h00230155;
         945:    rdata = 32'h4501000a;
         946:    rdata = 32'h446240f2;
         947:    rdata = 32'h494244d2;
         948:    rdata = 32'h4a2249b2;
         949:    rdata = 32'h61054a92;
         950:    rdata = 32'h04058082;
         951:    rdata = 32'h4505bfc9;
         952:    rdata = 32'h451cb7e5;
         953:    rdata = 32'h00b78023;
         954:    rdata = 32'h439c415c;
         955:    rdata = 32'h4817d793;
         956:    rdata = 32'h8082ffe5;
         957:    rdata = 32'hc4221141;
         958:    rdata = 32'hc606c226;
         959:    rdata = 32'h842e84aa;
         960:    rdata = 32'h00044583;
         961:    rdata = 32'h04058526;
         962:    rdata = 32'h47833fe9;
         963:    rdata = 32'hfbedfff4;
         964:    rdata = 32'h442240b2;
         965:    rdata = 32'h01414492;
         966:    rdata = 32'h415c8082;
         967:    rdata = 32'h89054388;
         968:    rdata = 32'hc10c8082;
         969:    rdata = 32'h8082c150;
         970:    rdata = 32'h99f14108;
         971:    rdata = 32'h8082952e;
         972:    rdata = 32'h80824148;
         973:    rdata = 32'h00a5c7b3;
         974:    rdata = 32'h0037f793;
         975:    rdata = 32'h00c508b3;
         976:    rdata = 32'h06079263;
         977:    rdata = 32'h00300793;
         978:    rdata = 32'h04c7fe63;
         979:    rdata = 32'h00357793;
         980:    rdata = 32'h00050713;
         981:    rdata = 32'h06079863;
         982:    rdata = 32'hffc8f613;
         983:    rdata = 32'hfe060793;
         984:    rdata = 32'h08f76c63;
         985:    rdata = 32'h02c77c63;
         986:    rdata = 32'h00058693;
         987:    rdata = 32'h00070793;
         988:    rdata = 32'h0006a803;
         989:    rdata = 32'h00478793;
         990:    rdata = 32'h00468693;
         991:    rdata = 32'hff07ae23;
         992:    rdata = 32'hfec7e8e3;
         993:    rdata = 32'hfff60793;
         994:    rdata = 32'h40e787b3;
         995:    rdata = 32'hffc7f793;
         996:    rdata = 32'h00478793;
         997:    rdata = 32'h00f70733;
         998:    rdata = 32'h00f585b3;
         999:    rdata = 32'h01176863;
        1000:    rdata = 32'h00008067;
        1001:    rdata = 32'h00050713;
        1002:    rdata = 32'hff157ce3;
        1003:    rdata = 32'h0005c783;
        1004:    rdata = 32'h00170713;
        1005:    rdata = 32'h00158593;
        1006:    rdata = 32'hfef70fa3;
        1007:    rdata = 32'hff1768e3;
        1008:    rdata = 32'h00008067;
        1009:    rdata = 32'h0005c683;
        1010:    rdata = 32'h00170713;
        1011:    rdata = 32'h00377793;
        1012:    rdata = 32'hfed70fa3;
        1013:    rdata = 32'h00158593;
        1014:    rdata = 32'hf80780e3;
        1015:    rdata = 32'h0005c683;
        1016:    rdata = 32'h00170713;
        1017:    rdata = 32'h00377793;
        1018:    rdata = 32'hfed70fa3;
        1019:    rdata = 32'h00158593;
        1020:    rdata = 32'hfc079ae3;
        1021:    rdata = 32'hf65ff06f;
        1022:    rdata = 32'h0045a683;
        1023:    rdata = 32'h0005a283;
        1024:    rdata = 32'h0085af83;
        1025:    rdata = 32'h00c5af03;
        1026:    rdata = 32'h0105ae83;
        1027:    rdata = 32'h0145ae03;
        1028:    rdata = 32'h0185a303;
        1029:    rdata = 32'h01c5a803;
        1030:    rdata = 32'h00d72223;
        1031:    rdata = 32'h0205a683;
        1032:    rdata = 32'h00572023;
        1033:    rdata = 32'h01f72423;
        1034:    rdata = 32'h01e72623;
        1035:    rdata = 32'h01d72823;
        1036:    rdata = 32'h01c72a23;
        1037:    rdata = 32'h00672c23;
        1038:    rdata = 32'h01072e23;
        1039:    rdata = 32'h02d72023;
        1040:    rdata = 32'h02470713;
        1041:    rdata = 32'h02458593;
        1042:    rdata = 32'hfaf768e3;
        1043:    rdata = 32'hf19ff06f;
        1044:    rdata = 32'h00f00313;
        1045:    rdata = 32'h00050713;
        1046:    rdata = 32'h02c37e63;
        1047:    rdata = 32'h00f77793;
        1048:    rdata = 32'h0a079063;
        1049:    rdata = 32'h08059263;
        1050:    rdata = 32'hff067693;
        1051:    rdata = 32'h00f67613;
        1052:    rdata = 32'h00e686b3;
        1053:    rdata = 32'h00b72023;
        1054:    rdata = 32'h00b72223;
        1055:    rdata = 32'h00b72423;
        1056:    rdata = 32'h00b72623;
        1057:    rdata = 32'h01070713;
        1058:    rdata = 32'hfed766e3;
        1059:    rdata = 32'h00061463;
        1060:    rdata = 32'h00008067;
        1061:    rdata = 32'h40c306b3;
        1062:    rdata = 32'h00269693;
        1063:    rdata = 32'h00000297;
        1064:    rdata = 32'h005686b3;
        1065:    rdata = 32'h00c68067;
        1066:    rdata = 32'h00b70723;
        1067:    rdata = 32'h00b706a3;
        1068:    rdata = 32'h00b70623;
        1069:    rdata = 32'h00b705a3;
        1070:    rdata = 32'h00b70523;
        1071:    rdata = 32'h00b704a3;
        1072:    rdata = 32'h00b70423;
        1073:    rdata = 32'h00b703a3;
        1074:    rdata = 32'h00b70323;
        1075:    rdata = 32'h00b702a3;
        1076:    rdata = 32'h00b70223;
        1077:    rdata = 32'h00b701a3;
        1078:    rdata = 32'h00b70123;
        1079:    rdata = 32'h00b700a3;
        1080:    rdata = 32'h00b70023;
        1081:    rdata = 32'h00008067;
        1082:    rdata = 32'h0ff5f593;
        1083:    rdata = 32'h00859693;
        1084:    rdata = 32'h00d5e5b3;
        1085:    rdata = 32'h01059693;
        1086:    rdata = 32'h00d5e5b3;
        1087:    rdata = 32'hf6dff06f;
        1088:    rdata = 32'h00279693;
        1089:    rdata = 32'h00000297;
        1090:    rdata = 32'h005686b3;
        1091:    rdata = 32'h00008293;
        1092:    rdata = 32'hfa0680e7;
        1093:    rdata = 32'h00028093;
        1094:    rdata = 32'hff078793;
        1095:    rdata = 32'h40f70733;
        1096:    rdata = 32'h00f60633;
        1097:    rdata = 32'hf6c378e3;
        1098:    rdata = 32'hf3dff06f;
        1099:    rdata = 32'h00b56733;
        1100:    rdata = 32'hfff00393;
        1101:    rdata = 32'h00377713;
        1102:    rdata = 32'h10071063;
        1103:    rdata = 32'h7f7f87b7;
        1104:    rdata = 32'hf7f78793;
        1105:    rdata = 32'h00052603;
        1106:    rdata = 32'h0005a683;
        1107:    rdata = 32'h00f672b3;
        1108:    rdata = 32'h00f66333;
        1109:    rdata = 32'h00f282b3;
        1110:    rdata = 32'h0062e2b3;
        1111:    rdata = 32'h10729263;
        1112:    rdata = 32'h08d61663;
        1113:    rdata = 32'h00452603;
        1114:    rdata = 32'h0045a683;
        1115:    rdata = 32'h00f672b3;
        1116:    rdata = 32'h00f66333;
        1117:    rdata = 32'h00f282b3;
        1118:    rdata = 32'h0062e2b3;
        1119:    rdata = 32'h0c729e63;
        1120:    rdata = 32'h06d61663;
        1121:    rdata = 32'h00852603;
        1122:    rdata = 32'h0085a683;
        1123:    rdata = 32'h00f672b3;
        1124:    rdata = 32'h00f66333;
        1125:    rdata = 32'h00f282b3;
        1126:    rdata = 32'h0062e2b3;
        1127:    rdata = 32'h0c729863;
        1128:    rdata = 32'h04d61663;
        1129:    rdata = 32'h00c52603;
        1130:    rdata = 32'h00c5a683;
        1131:    rdata = 32'h00f672b3;
        1132:    rdata = 32'h00f66333;
        1133:    rdata = 32'h00f282b3;
        1134:    rdata = 32'h0062e2b3;
        1135:    rdata = 32'h0c729263;
        1136:    rdata = 32'h02d61663;
        1137:    rdata = 32'h01052603;
        1138:    rdata = 32'h0105a683;
        1139:    rdata = 32'h00f672b3;
        1140:    rdata = 32'h00f66333;
        1141:    rdata = 32'h00f282b3;
        1142:    rdata = 32'h0062e2b3;
        1143:    rdata = 32'h0a729c63;
        1144:    rdata = 32'h01450513;
        1145:    rdata = 32'h01458593;
        1146:    rdata = 32'hf4d60ee3;
        1147:    rdata = 32'h01061713;
        1148:    rdata = 32'h01069793;
        1149:    rdata = 32'h00f71e63;
        1150:    rdata = 32'h01065713;
        1151:    rdata = 32'h0106d793;
        1152:    rdata = 32'h40f70533;
        1153:    rdata = 32'h0ff57593;
        1154:    rdata = 32'h02059063;
        1155:    rdata = 32'h00008067;
        1156:    rdata = 32'h01075713;
        1157:    rdata = 32'h0107d793;
        1158:    rdata = 32'h40f70533;
        1159:    rdata = 32'h0ff57593;
        1160:    rdata = 32'h00059463;
        1161:    rdata = 32'h00008067;
        1162:    rdata = 32'h0ff77713;
        1163:    rdata = 32'h0ff7f793;
        1164:    rdata = 32'h40f70533;
        1165:    rdata = 32'h00008067;
        1166:    rdata = 32'h00054603;
        1167:    rdata = 32'h0005c683;
        1168:    rdata = 32'h00150513;
        1169:    rdata = 32'h00158593;
        1170:    rdata = 32'h00d61463;
        1171:    rdata = 32'hfe0616e3;
        1172:    rdata = 32'h40d60533;
        1173:    rdata = 32'h00008067;
        1174:    rdata = 32'h00450513;
        1175:    rdata = 32'h00458593;
        1176:    rdata = 32'hfcd61ce3;
        1177:    rdata = 32'h00000513;
        1178:    rdata = 32'h00008067;
        1179:    rdata = 32'h00850513;
        1180:    rdata = 32'h00858593;
        1181:    rdata = 32'hfcd612e3;
        1182:    rdata = 32'h00000513;
        1183:    rdata = 32'h00008067;
        1184:    rdata = 32'h00c50513;
        1185:    rdata = 32'h00c58593;
        1186:    rdata = 32'hfad618e3;
        1187:    rdata = 32'h00000513;
        1188:    rdata = 32'h00008067;
        1189:    rdata = 32'h01050513;
        1190:    rdata = 32'h01058593;
        1191:    rdata = 32'hf8d61ee3;
        1192:    rdata = 32'h00000513;
        1193:    rdata = 32'h00008067;
        1194:    rdata = 32'h05971101;
        1195:    rdata = 32'h85930000;
        1196:    rdata = 32'hf5171165;
        1197:    rdata = 32'h0513000e;
        1198:    rdata = 32'hce06d9a5;
        1199:    rdata = 32'h00683925;
        1200:    rdata = 32'h854ff0ef;
        1201:    rdata = 32'h450140f2;
        1202:    rdata = 32'h80826105;
        1203:    rdata = 32'h010005b7;
        1204:    rdata = 32'h000ef517;
        1205:    rdata = 32'hd3050513;
        1206:    rdata = 32'h95dff06f;
        1207:    rdata = 32'h010105b7;
        1208:    rdata = 32'h000ef517;
        1209:    rdata = 32'hd4050513;
        1210:    rdata = 32'h9e5ff06f;
        1211:    rdata = 32'h010025b7;
        1212:    rdata = 32'h000ef517;
        1213:    rdata = 32'hd5c50513;
        1214:    rdata = 32'hf797beb9;
        1215:    rdata = 32'h8793000e;
        1216:    rdata = 32'h6741d727;
        1217:    rdata = 32'h6711c398;
        1218:    rdata = 32'h8082c3d8;
        1219:    rdata = 32'h00000000;
        1220:    rdata = 32'h00000000;
        1221:    rdata = 32'h00000000;
        1222:    rdata = 32'h00000000;
        1223:    rdata = 32'h000112cc;
        1224:    rdata = 32'h000112dc;
        1225:    rdata = 32'h000112ec;
        1226:    rdata = 32'h000112fa;
        1227:    rdata = 32'hfffff026;
        1228:    rdata = 32'hfffff02c;
        1229:    rdata = 32'hfffff032;
        1230:    rdata = 32'hfffff038;
        1231:    rdata = 32'hfffff03e;
        1232:    rdata = 32'h0002c000;
        1233:    rdata = 32'h0003c000;
        1234:    rdata = 32'hc00002c0;
        1235:    rdata = 32'h02c00003;
        1236:    rdata = 32'h0003c000;
        1237:    rdata = 32'hc00002c0;
        1238:    rdata = 32'h02c00003;
        1239:    rdata = 32'h0003c000;
        1240:    rdata = 32'hc00002c0;
        1241:    rdata = 32'h02c00003;
        1242:    rdata = 32'h0003c000;
        1243:    rdata = 32'hc00002c0;
        1244:    rdata = 32'h02c00003;
        1245:    rdata = 32'h0003c000;
        1246:    rdata = 32'hc00002c0;
        1247:    rdata = 32'h02c00003;
        1248:    rdata = 32'h0003c000;
        1249:    rdata = 32'hc00002c0;
        1250:    rdata = 32'h02c00003;
        1251:    rdata = 32'h0003c000;
        1252:    rdata = 32'hc00002c0;
        1253:    rdata = 32'h02c00003;
        1254:    rdata = 32'h0003c000;
        1255:    rdata = 32'hc00002c0;
        1256:    rdata = 32'h02c00003;
        1257:    rdata = 32'h00042000;
        1258:    rdata = 32'h0020c000;
        1259:    rdata = 32'h200000c0;
        1260:    rdata = 32'h00000000;
        1261:    rdata = 32'h0008c000;
        1262:    rdata = 32'h200000c0;
        1263:    rdata = 32'h00000000;
        1264:    rdata = 32'h6c707061;
        1265:    rdata = 32'h74616369;
        1266:    rdata = 32'h206e6f69;
        1267:    rdata = 32'h72617473;
        1268:    rdata = 32'h0a646574;
        1269:    rdata = 32'h00000000;
        1270:    rdata = 32'h0000203e;
        1271:    rdata = 32'h706c6568;
        1272:    rdata = 32'h20202020;
        1273:    rdata = 32'h20202020;
        1274:    rdata = 32'h20202020;
        1275:    rdata = 32'h70202d20;
        1276:    rdata = 32'h746e6972;
        1277:    rdata = 32'h69687420;
        1278:    rdata = 32'h656d2073;
        1279:    rdata = 32'h67617373;
        1280:    rdata = 32'h65730a65;
        1281:    rdata = 32'h656c5f74;
        1282:    rdata = 32'h20202064;
        1283:    rdata = 32'h20202020;
        1284:    rdata = 32'h2d202020;
        1285:    rdata = 32'h74657320;
        1286:    rdata = 32'h64656c20;
        1287:    rdata = 32'h6165720a;
        1288:    rdata = 32'h616d5f64;
        1289:    rdata = 32'h78697274;
        1290:    rdata = 32'h20202020;
        1291:    rdata = 32'h202d2020;
        1292:    rdata = 32'h64616572;
        1293:    rdata = 32'h74616d20;
        1294:    rdata = 32'h0a786972;
        1295:    rdata = 32'h696c6163;
        1296:    rdata = 32'h74617262;
        1297:    rdata = 32'h616d5f65;
        1298:    rdata = 32'h78697274;
        1299:    rdata = 32'h63202d20;
        1300:    rdata = 32'h62696c61;
        1301:    rdata = 32'h65746172;
        1302:    rdata = 32'h78697020;
        1303:    rdata = 32'h20736c65;
        1304:    rdata = 32'h7366666f;
        1305:    rdata = 32'h0a737465;
        1306:    rdata = 32'h00000000;
        1307:    rdata = 32'h006e6970;
        1308:    rdata = 32'h74617473;
        1309:    rdata = 32'h00000065;
        1310:    rdata = 32'h64616572;
        1311:    rdata = 32'h5f74756f;
        1312:    rdata = 32'h656d6974;
        1313:    rdata = 32'h00000000;
        1314:    rdata = 32'h7366666f;
        1315:    rdata = 32'h63207465;
        1316:    rdata = 32'h62696c61;
        1317:    rdata = 32'h69746172;
        1318:    rdata = 32'h64206e6f;
        1319:    rdata = 32'h0a656e6f;
        1320:    rdata = 32'h00000000;
        1321:    rdata = 32'h696c6163;
        1322:    rdata = 32'h74617262;
        1323:    rdata = 32'h5f6e6f69;
        1324:    rdata = 32'h656d6974;
        1325:    rdata = 32'h00000000;
        1326:    rdata = 32'h65726e75;
        1327:    rdata = 32'h6e676f63;
        1328:    rdata = 32'h64657a69;
        1329:    rdata = 32'h6d6f6320;
        1330:    rdata = 32'h646e616d;
        1331:    rdata = 32'h0000000a;
        1332:    rdata = 32'h706c6568;
        1333:    rdata = 32'h00000000;
        1334:    rdata = 32'h5f746573;
        1335:    rdata = 32'h0064656c;
        1336:    rdata = 32'h64616572;
        1337:    rdata = 32'h74616d5f;
        1338:    rdata = 32'h00786972;
        1339:    rdata = 32'h696c6163;
        1340:    rdata = 32'h74617262;
        1341:    rdata = 32'h616d5f65;
        1342:    rdata = 32'h78697274;
        1343:    rdata = 32'h00000000;
        1344:    rdata = 32'h0000203a;
        1345:    rdata = 32'h00002820;
        1346:    rdata = 32'h00203a29;
        1347:    rdata = 32'h6f636e69;
        1348:    rdata = 32'h63657272;
        1349:    rdata = 32'h61762074;
        1350:    rdata = 32'h2e65756c;
        1351:    rdata = 32'h79727420;
        1352:    rdata = 32'h61676120;
        1353:    rdata = 32'h000a6e69;
        default: rdata = 32'h00000000;
    endcase
end
endmodule
