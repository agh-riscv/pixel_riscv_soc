/**
 * Copyright (C) 2020  AGH University of Science and Technology
 *
 * This program is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with this program.  If not, see <https://www.gnu.org/licenses/>.
 */

module boot_rom (
    input logic          clk,
    input logic          rst_n,
    ibex_data_bus.slave  data_bus,
    ibex_instr_bus.slave instr_bus
);


/**
 * Local variables and signals
 */

typedef enum logic [1:0] {
    IDLE,
    DATA_READOUT,
    INSTR_READOUT
} state_t;


/**
 * Local variables and signals
 */

state_t      state, state_nxt;
logic [31:0] addr, rdata;


/**
 * Signals assignments
 */

assign data_bus.rdata_intg = 7'b0;
assign data_bus.err = 1'b0;

assign instr_bus.rdata_intg = 7'b0;
assign instr_bus.err = 1'b0;


/**
 * Submodules placement
 */

boot_mem u_boot_mem (
    .rdata,
    .addr
);


/**
 * Module internal logic
 */

always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n)
        state <= IDLE;
    else
        state <= state_nxt;
end

always_comb begin
    state_nxt = state;

    case (state)
    IDLE: begin
        if (data_bus.req)
            state_nxt = DATA_READOUT;
        else if (instr_bus.req)
            state_nxt = INSTR_READOUT;
    end
    DATA_READOUT,
    INSTR_READOUT: begin
        state_nxt = IDLE;
    end
    endcase
end

always_comb begin
    data_bus.gnt = 1'b0;
    instr_bus.gnt = 1'b0;

    case (state)
    IDLE: begin
        if (data_bus.req)
            data_bus.gnt = 1'b1;
        else if (instr_bus.req)
            instr_bus.gnt = 1'b1;
    end
    DATA_READOUT,
    INSTR_READOUT: ;
    endcase
end

always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        addr <= 32'b0;
    end else begin
        case (state)
        IDLE: begin
            if (data_bus.req)
                addr <= data_bus.addr;
            else if (instr_bus.req)
                addr <= instr_bus.addr;
        end
        DATA_READOUT,
        INSTR_READOUT: ;
        endcase
    end
end

always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        data_bus.rvalid <= 1'b0;
        data_bus.rdata <= 32'b0;
        instr_bus.rvalid <= 1'b0;
        instr_bus.rdata <= 32'b0;
    end else begin
        case (state)
        IDLE: begin
            data_bus.rvalid <= 1'b0;
            instr_bus.rvalid <= 1'b0;
        end
        DATA_READOUT: begin
            data_bus.rvalid <= 1'b1;
            data_bus.rdata <= rdata;
        end
        INSTR_READOUT: begin
            instr_bus.rvalid <= 1'b1;
            instr_bus.rdata <= rdata;
        end
        endcase
    end
end

endmodule
